localparam  MAJOR_VERSION='h0;
localparam  MINOR_VERSION='h5;
localparam  REVISION_NUM='h3;
localparam  DEBUG_REVISION='h0;
localparam  FH_MODE='h1;
localparam  NUM_ETH_CORES='h2;
localparam  FDD_SUPPORTED='h0;
localparam  TDD_SUPPORTED='h1;
localparam  MAX_SUPPORTED_ANTENNAS='h8;
localparam  MAX_SUPPORTED_CARRIERS='h2;
localparam  MAX_PRECISION='h16;
localparam  CAR0_LTE_SUPPORTED='h0;
localparam  CAR1_LTE_SUPPORTED='h0;
localparam  CAR0_5G_SUPPORTED='h1;
localparam  CAR1_5G_SUPPORTED='h1;
localparam  NUMEROLOGY0_SUPPORTED='h0;
localparam  NUMEROLOGY1_SUPPORTED='h1;
localparam  NUMEROLOGY2_SUPPORTED='h0;
localparam  EXTENDED_CP_SUPPORTED='h0;
localparam  SEC_TYPE0_SUPPORTED='h1;
localparam  SEC_TYPE1_SUPPORTED='h1;
localparam  SEC_TYPE3_SUPPORTED='h1;
localparam  CAR0_PRACH_LTE_FORMAT0_SUPPORTED='h0;
localparam  CAR0_PRACH_LTE_FORMAT1_SUPPORTED='h0;
localparam  CAR0_PRACH_LTE_FORMAT2_SUPPORTED='h0;
localparam  CAR0_PRACH_LTE_FORMAT3_SUPPORTED='h0;
localparam  CAR0_PRACH_LTE_FORMAT4_SUPPORTED='h0;
localparam  CAR1_PRACH_LTE_FORMAT0_SUPPORTED='h0;
localparam  CAR1_PRACH_LTE_FORMAT1_SUPPORTED='h0;
localparam  CAR1_PRACH_LTE_FORMAT2_SUPPORTED='h0;
localparam  CAR1_PRACH_LTE_FORMAT3_SUPPORTED='h0;
localparam  CAR1_PRACH_LTE_FORMAT4_SUPPORTED='h0;
localparam  CAR0_PRACH_5G_FORMAT0_SUPPORTED='h1;
localparam  CAR0_PRACH_5G_FORMAT1_SUPPORTED='h0;
localparam  CAR0_PRACH_5G_FORMAT2_SUPPORTED='h0;
localparam  CAR0_PRACH_5G_FORMAT3_SUPPORTED='h0;
localparam  CAR1_PRACH_5G_FORMAT0_SUPPORTED='h1;
localparam  CAR1_PRACH_5G_FORMAT1_SUPPORTED='h0;
localparam  CAR1_PRACH_5G_FORMAT2_SUPPORTED='h0;
localparam  CAR1_PRACH_5G_FORMAT3_SUPPORTED='h0;
localparam  CAR0_BW_5MHZ_SUPPORTED='h0;
localparam  CAR0_BW_10MHZ_SUPPORTED='h0;
localparam  CAR0_BW_15MHZ_SUPPORTED='h0;
localparam  CAR0_BW_20MHZ_SUPPORTED='h0;
localparam  CAR0_BW_40MHZ_SUPPORTED='h0;
localparam  CAR0_BW_60MHZ_SUPPORTED='h0;
localparam  CAR0_BW_80MHZ_SUPPORTED='h0;
localparam  CAR0_BW_100MHZ_SUPPORTED='h1;
localparam  CAR1_BW_5MHZ_SUPPORTED='h0;
localparam  CAR1_BW_10MHZ_SUPPORTED='h0;
localparam  CAR1_BW_15MHZ_SUPPORTED='h0;
localparam  CAR1_BW_20MHZ_SUPPORTED='h0;
localparam  CAR1_BW_40MHZ_SUPPORTED='h0;
localparam  CAR1_BW_60MHZ_SUPPORTED='h0;
localparam  CAR1_BW_80MHZ_SUPPORTED='h0;
localparam  CAR1_BW_100MHZ_SUPPORTED='h1;
localparam  T2A_MIN_UP_NS_100MHZ='h1C138;
localparam  T2A_MIN_UP_NS_80MHZ='h1C138;
localparam  T2A_MIN_UP_NS_60MHZ='h1C138;
localparam  T2A_MIN_UP_NS_40MHZ='h1C138;
localparam  T2A_MIN_UP_NS_20MHZ='h1C138;
localparam  T2A_MIN_UP_NS_15MHZ='h1C138;
localparam  T2A_MIN_UP_NS_10MHZ='h1D293;
localparam  T2A_MIN_UP_NS_5MHZ='h1F377;
localparam  TUP_RECEPTION_WINDOW_DL_NS='h72038;
localparam  TCP_RECEPTION_WINDOW_DL_NS='h48440;
localparam  TCP_ADV_DL_NS='h1D4C0;
localparam  TA3_MIN_UP_NS_100MHZ='h1D79C;
localparam  TA3_MIN_UP_NS_80MHZ='h1D79C;
localparam  TA3_MIN_UP_NS_60MHZ='h1D79C;
localparam  TA3_MIN_UP_NS_40MHZ='h1D79C;
localparam  TA3_MIN_UP_NS_20MHZ='h1D79C;
localparam  TA3_MIN_UP_NS_15MHZ='h1D79C;
localparam  TA3_MIN_UP_NS_10MHZ='h21ABF;
localparam  TA3_MIN_UP_NS_5MHZ='h1E908;
localparam  TA3_MIN_UP_PRACH_NS_100MHZ='h15DD2;
localparam  TA3_MIN_UP_PRACH_NS_80MHZ='h15DD2;
localparam  TA3_MIN_UP_PRACH_NS_60MHZ='h15DD2;
localparam  TA3_MIN_UP_PRACH_NS_40MHZ='h15DD2;
localparam  TA3_MIN_UP_PRACH_NS_20MHZ='h15DD2;
localparam  TA3_MIN_UP_PRACH_NS_15MHZ='h15DD2;
localparam  TA3_MIN_UP_PRACH_NS_10MHZ='h169DE;
localparam  TA3_MIN_UP_PRACH_NS_5MHZ='h19A4F;
localparam  TUP_TRANSMISSION_WINDOW_UL_NS='h7918;
localparam  T2A_MIN_CP_UL_NS='h0;
localparam  TCP_RECEPTION_WINDOW_UL_NS='h81A38;
localparam  DL_FRM_MRKR_TIME_ADVANCE_100MHZ='h1AAC8;
localparam  DL_FRM_MRKR_TIME_ADVANCE_80MHZ='h1AAC8;
localparam  DL_FRM_MRKR_TIME_ADVANCE_60MHZ='h1AAC8;
localparam  DL_FRM_MRKR_TIME_ADVANCE_40MHZ='h1AAC8;
localparam  DL_FRM_MRKR_TIME_ADVANCE_20MHZ='h1AAC8;
localparam  DL_FRM_MRKR_TIME_ADVANCE_15MHZ='h1AAC8;
localparam  DL_FRM_MRKR_TIME_ADVANCE_10MHZ='h1BC6C;
localparam  DL_FRM_MRKR_TIME_ADVANCE_5MHZ='h1DD4F;
localparam  UL_FRM_MRKR_TIME_DELAY_100MHZ='hEDC;
localparam  UL_FRM_MRKR_TIME_DELAY_80MHZ='hEDC;
localparam  UL_FRM_MRKR_TIME_DELAY_60MHZ='hEDC;
localparam  UL_FRM_MRKR_TIME_DELAY_40MHZ='hEDC;
localparam  UL_FRM_MRKR_TIME_DELAY_20MHZ='hEDC;
localparam  UL_FRM_MRKR_TIME_DELAY_15MHZ='hEDC;
localparam  UL_FRM_MRKR_TIME_DELAY_10MHZ='h1B62;
localparam  UL_FRM_MRKR_TIME_DELAY_5MHZ='h333A;
localparam  PRACH_FRM_MRKR_TIME_DELAY_100MHZ='h12CF0;
localparam  PRACH_FRM_MRKR_TIME_DELAY_80MHZ='h12CF0;
localparam  PRACH_FRM_MRKR_TIME_DELAY_60MHZ='h12CF0;
localparam  PRACH_FRM_MRKR_TIME_DELAY_40MHZ='h12CF0;
localparam  PRACH_FRM_MRKR_TIME_DELAY_20MHZ='h12CF0;
localparam  PRACH_FRM_MRKR_TIME_DELAY_15MHZ='h12CF0;
localparam  PRACH_FRM_MRKR_TIME_DELAY_10MHZ='h138FC;
localparam  PRACH_FRM_MRKR_TIME_DELAY_5MHZ='h1696D;
localparam  TSSI_SAMPLES_PER_15P36_TIC='h20;
localparam  TSSI_ACCUM_TRUNCATED_BITS='h19;
localparam  WRSSI_SAMPLES_PER_15P36_TIC='h20;
localparam  WRSSI_ACCUM_TRUNCATED_BITS='h19;
localparam  RSSI_SAMPLES_PER_15P36_TIC_20M='h2;
localparam  RSSI_ACCUM_TRUNCATED_BITS='h19;
localparam  CFR_SAMPLE_PERIOD_PS='h7F2;
localparam  PATH_DELAY_SAMPLE_PERIOD_PS='h1FCA;
localparam  DL_TIME_DELAY_BYPASS='h0;
localparam  UL_TIME_DELAY_BYPASS='h0;

`define RSP_S2_DMA_SECT_BASE_ADDR                                   'h0
`define RSP_S2_DMA_CSR_REG_CSR0_BASE_ADDR                           'h0
`define RSP_S2_DMA_CSR_REG_CSR0_END_ADDR                            'h3ff
`define RSP_S2_DMA_CSR_REG_CSR1_BASE_ADDR                           'h400
`define RSP_S2_DMA_CSR_REG_CSR1_END_ADDR                            'h7ff
`define RSP_S2_DMA_CSR_REG_CSR2_BASE_ADDR                           'h800
`define RSP_S2_DMA_CSR_REG_CSR2_END_ADDR                            'hbff
`define RSP_S2_DMA_CSR_REG_CSR3_BASE_ADDR                           'hc00
`define RSP_S2_DMA_CSR_REG_CSR3_END_ADDR                            'hfff
`define RSP_S2_DMA_GLB_REG_BASE_ADDR                                'h1000
`define RSP_S2_DMA_GLB_REG_END_ADDR                                 'h13ff


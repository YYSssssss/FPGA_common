`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
ph4fbHMLdHMt9t3rD6l++tYcXEMDkmgkdD4mqYPn5Ze35RUC0m4kgOryQJwBCU+MP5iDaTYYRV5g
4SWI0DkcpQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
p3MoKO2wTFS+7WBVYUX0FOz9xBvTflfGDUU+W62MMVogCsaiuXr6A5NK3Y6MmhqxZGkElHofu+sf
FxtOG7CavHmqJtttKJfk9jzLq6DGYjvPrhDLfonBFJ7+qWzop9HKJW3IAIyPBrOX57C3hWf5T658
fwIou8Pk1CYK1P9flps=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
En2AK/Wgqk2oLRY5SjEfmbRdpDPJJgf7r2ZCEonj0CmHo3+r7CvDsdWlpsV2KlSuYhtpeX+vuwVn
2qQMzPyxnS2YcpmizlDVWOvi0zV4dRjj7r4CCVcKb/9Wg04VnnxoLgFbyxpZ6n8uA0eWuwHzC8Yl
Z8dzu6JMOi6EO/x4ZcIiI8MJiyOboyVzyx7V+ja+eS87qowm7tAroCckmNEYOvARBFQmT1AtIHSy
dyOlUEbZIpp0vqV6OpKK6Rr8wiLfCKJqkomGF40yx5rsJ+8bNlgg6udeFS0x41q6T3//RHoERzWI
FTeKY1UlAiB+ytKEUUtCnwQD1iwFGQgfJ0h2Kw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fPd069tEZZz5v2NgXzRiuqS2lAEPLCdDDXFukVTw71UsqqbYLfeXFaPaXoa02TcQZrydmutcrtlR
J/26u3DYVea+zJKTBjcHqbaopWcTiU18NJgULOCQOWFJqPgyEhxXpIvd2ETbgpM+ifWoInP8dUlD
8GhUSqmk3Zup15GmhfmNSPFeHlAaXNEYCxS64VLPPqO270tzzX2ffgkpfjih3XEBOEWV2/fRMEIU
3Np97+pUw2m+IJwt/HQ4PJVtGygekdul8yF751pcjPuaryGDM85zzRgGFhGSovp6sBFcDSlu3Jvt
adzhldYd0ezTTk4relN5Br4pkujkM6OY4X90wg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
tR7PxLcMjSI9wwUgk9tTHdcY8Uwia2NXW5kaLvO9gswxN1GtL9GSPgbb5zr+sTnp/S+LKTI+02KI
TMB2geQgK1pZkvdk0+Ol3vq6Tk3Zk42Qe74Vf2ZvuojvmkV2QKZFg/aa2tb5O17kne5a1IXrg8l5
z6Yi8tPHSXCNwciJWpk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Bds0en+2c8yztwhHVpMedOFRj8NmE/EEWnfaOlQDyHm80o1CcC4cZHg54ZpJfMa9/U+YW6bNpsqS
FhcQ+qEiE6QQJpUFJJDqKhpO5QotCv5d1x0qrjaitJ2226PAPA9tN8Z/ZVce7wJ2S3dwf9yv+8dO
rbJQQd2+lF8shy5foQRER8hcOnAeL0MibzMiJVU86M0mN3Iy0EBiQ53foAu5et5iMNly+0Z9/L1h
C7LP+1MRwZ+VA/mHmo+cKOnpQvLRRhGLaMCOfV7WF96dPXwZ3Z0TmQJx7RSddqeV9LftOvrNpRPm
aZmc0GNJbK+RYV604McyE2SwMEOkx3LMghALCg==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
alO/bSTeEnbogP4KcCzgjgW1pQWnX9Bgzz3D9ibL100OPGDpXUyCgBBmGhN1F+GR4iwTbtF8aSP6
YKMJKr+0QUueXQWwattLlV/7yK4r+c6cmCm0MCVhnSiJHVen61GwWEUTqOKfd994wP7ZJbNdNk5n
0JP5kG6akdfavqt2saV1wC9SH3QphpL2qBB5dgec2Wn9Z6tERWnKrNCXCbntKuofu8/rom6f7/AW
I8Dd6ms+fvD2PL25Z6FKZSFzf/u0leeiQUpvB2Mhe5gCIymdEICsjronnhzSfBZmmx1qDmPXHc7L
uU6kVDl3MNUB3mCc4AvJCIdEErJ1cH9EPBaf0g==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KCBkW2omby+FZy53+sB2qtEp1Oa8tM9yMQWpQaEh4yvplMjPiDdlXmiSm4hbpZLfNX3IaW8TSza0
oFxVjuH7/T+WzbOgY/r6i1SoZuE8NtexB7fAymGCfsDcRvuRFBDUt9jmkNxiuuHL4aVNl5gU67Jp
sBl16ERKxQGL94PtR3xNLEYFXxkSYXrIciqnbXyU9KqS0axlAHXIEOK7mm/hsRsRj06sh0uSf7AO
DH002lKncjh5xlS+ad/B3fX+vaA1r0RdEf4gN1nATKsquH+Ezcunc13CjIsU6WmSMjDcr2wjM1+V
x5raLGvn37SSxXKBZRGMYMEnl+M0CNQMgcbI8A==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OKpvCZ5EyJbwgo77eKHb/YSI/lADZw0WqLSeEIH3GOBl5NeXzWp8RRMTLyWMYeG4JehSE9jn1nM8
FPbheCZKwZBAFYyZ4rgE8YGf/ykvuflSJm2uXugw2Cn/Zr84QaKZ1e+OCPoqJXO7IVVpzu/1/c5e
t199mzUJEQbmVnBy09AgqYRqBFElANrfIvkBxa5u2kh6Q3gKrFXeXiFGDdDoW9xvShdZClFR0eSg
MDl3FGGLguyTSZWrFdkpgryN6kpruoRCKFntoicEsRcte8ecJZhgcNsC2XMgZHGFHn4i+mQSQkM+
f05kNS9z3oa05gupkS5T7eunOYwPfeAooMVZHQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 82320)
`pragma protect data_block
RfYxomztYJaIWoKVoB+VWmjoZKD6Wcz15a8w4wbJSTe8VXFH4wvluS0Hx+E5f3E4s0F7BQQnyyY+
XM8gR5uM/UwPl3PgmJrybSPkRpG0xEEFoaH4HozwasS/farGbgI8SSaKyRhkh8N/EGG7GAp2pFOO
S7wmjc8KId0+GT35MOYyiR+BGntiTIS+PzrQz8wmQ3ANS2SfZTYZKdmqv0B8b9vzY4/WDmaXNKS6
7D82nCo9L7gCiH/oGBdWrh+vCfwrRg+k8ofI/EcQWT+7n3oVSV3k2IBe5qYtG29/nFiIFqC3BOmV
9dGUSYXBarJUe8RpRfhCV1n1JkGp5b6NM+YsUJMRA/et9EXVJRuZpj03QEZz6lLs6RvQxShDeGkm
BWMlYE5MmKHb0ePv5DAVrvO9K2mgr3Rs42FmtdoLbUsV5MJ9eKDwQUMQJASNVs4XNfNncMpLFG2e
z9jEKc/NVh8GOltYHWIepnt40MG5hQsfYUwf2Qk/pl4wA5qhoHYnQnn29KF4SD2jo/e6kWE3BRPr
WdChNUx6pjpvMEeh+6k1rAL0qh5E383k2qwxoraWonCa8O39IfoHG3a7drtgF+b1wuEzUAs1yaIg
BNCZ+KEYghKjKEgmdAhGwtqEq9sIMeisjpI1hl1k0DkIlISkmJBDgztN0l+qIsq0WfrmxMBZA7sl
Gz34dzEi2txEcSdia/cbKNHUSvVQftxsL7LBAAnw5jVtsbZsoIrhiY9+ja9seOg12mhqtL4wPNa9
gubc+zI7numm5WfPmvJ4ZV+k6ep431WOOF+G9m3RD6UK8czCBNyDUPNjjp1lORenBZM+Odx7zHJD
rRMwYIOijfjhdezqr45IyqcuZCUhttwOAgbLsav8445PVSc/R4n4gvrZb6dAOvYHFJdo0HjBWm6d
NsGcEx6bOgg0d0jNriSp7AnIggF/g4M30ACmZ1j0CJOA2TsE7E00DDg84n9qZDXq6iySHVpkNv02
No46vWOWKiFDyE6PwfYfQGx9wStpeDVQAAFhZ65CHLmcelKH1Dg73nSZT0Rsqmuncx9xMALgecZZ
wT1bewTNu1wlc/Tx8B23IoPu6ezGtmSH10qEFKyogNPxkvCdgCexT+SjLvo/YqsJYLPQ9n0LDczX
8/nAAZeaXaXuP1D2hZHQzGWg6lTKF1Z61b9Kli/XPaz+T5vOzqqMZje1xO0PR9BVO7QwpuI0TAfH
mGH2IoLbw/NoCddcqaH9ZWIEtBICoCqbuW3C9BETysPNblzgrWSm9GhgEDuk1VdiFTxSESBWllwS
RlDVMeyDdiYEpNwWY5K/HQdSL7DTe42wQp7mVSrXB61/xYp8bAFFsdJRnAvGTimoaRBwqqcE6r2X
//Jpm6MWdlQ/Km9C6OBLYuoNuuRtM52jqF4g89xWAPO+/4FrJA/eLKmue45UrdfCLTUejMbCdXGu
bx3S6zxRNgmJP+cPuz1g38fK+sWZH5UB9jutTvkdGJd/Z/OuNuK3yQxb5Z5AW6DQcy02jk0AVp6y
hqA81ihB/Ieb/9iGGZYHgOmoh04a2trg8mHWL9yhGNlWf1JeAxftux4GNhSBLoSncOljlfiGHAQq
xpL06dPcz/XEEWfP/KFBhK4ZMy4FlczbvEnUZOcyHz7DXEehbJ48aNh5RLTXUvDazL4McCuQ6StT
SPtj6uvLGiGfgo+FuJTWCrzfzEmLnYg9x0p77r3SmJF83+E72PBDk20gLeXDWVehBoYoAEo/zP88
cSFnkmrAqxa8gWWAMtr0bf373h6ilCM3pvPuxnbTamcSvn/+h8davtIRVyw+NVQINJgsARjrd8JL
qt/Yp2I8S1hX2igEKhmOTT/Cp2iJ0paKCe+In/M6VmN6Cgz9AY9g7z6Subf3WEc9pCK6E3peRHuR
GvKL6QSiqWySZlSHrN3nYDEbfRHh4INUZfvY1uHYy6uH3Bpuu8OoWQgI+qV6FzTCdvf3j73tQIYE
E8YSd78+0PDzmHrdRDxCscHU9qM+yQdhIBLMnCBMsnUC7AyBszdJO201ztejniwAWi4bHJpWEblN
WS2STaLTtsdtAztXUlKf3okPhup+8Qt9Oa1+/NaIxpu3hCdCAq1LPkvMv/zKMg4YwMlgmm6HVXEf
6LCgIn+X2c/8tvT7Y1RuClOae66NKE4pidz2xQqdDZn3625V+45X4b+bHw1I0RVqRyLbO5D6E0BK
EdpQbGWmE9DrSEBKL4UOufOHv9Fc0gclvbrMg8wyH3j1dN0TTJlz3mFM6mPcol/9kGKHIKJ5CDQ0
HY/6DEWfyrDNfTO/eAtMuzDM4jjq/cTmzYLyM/I5We2eH1ATB5Ke7cTbqq7yQbJFuqz0Zmhc4QmG
PvL0kuW5HSrXXQ6TUu4KUWqpTYUryJuUsw7QXESi/OjqV2NrA+vgL9lNEdrDuMV1V1t5jx6YkPGt
1pkgzgsTLOFG0uvM7AOaE7+Qgj39RDw0Kw8YEDJfKJUq+d/RPGKbdqX1OFQoFo3Vmg6WIQ2ptgO6
CkUtWL/EDBTPulB6sDJ6FgOsHtxKyIk/ZrtBDDGjolADpPQgylB2J6bXUVe1t3c/VN4GxwRE33wN
lsh4QU7c/SAr2S9XaAKLH7Sd6EGjbmNVwrOzjrL9EKuVosnQSwNEjkP4EusYzMscu3EZFjEXk+24
fzJbMWYGzSQvZXHU3WlqfFYbG4mQBeOKKw3X1k1a0GekP8iWEDKSaidpMo0rE8JFeCLUOsPxz5Bw
41bqp/XQvlFE5YjQQOh9sh4EMchbWJGbIhuKiQjHvfZv33t57StnY+FOLtSMvjPkGIk/tPdPfSmd
J6eDsTF4QSo2mkdzMirOHbEXrQMuebAkY2vZtA8++41PE5YsbLUwBUsiOO/e1iOu0vTC9RDnUHiz
cXGM6/l1TX3laXoIzARFrD9JuR76CP21WcMyVwJVe2//5ZMR4m8Dnf7UoD0l+EXP5VDf+1YjafKB
D3caE4YnXHSgraZ1C4eAo9X9M7Wy/qcL8UjSVMUwlqLpyt0JP9FSgid6HKiXndE2GLrTQ/5qMCsg
tWuRJTcZ1YczRlSxqlMrC65g65G2zNeSWQ//rJ1raJewSz8BL5Gcs2MouJG4ewsqbQyWUo2tsmxG
V/xM8aV8O4ENYXamhyXdfBXIgGt1NjD8wKgO3gIHoRaMn1YsdtuTofKyO/wKaItRNCuhxIYZyK9j
fNDHVzIAeBgz3H+R4DTLbF1QqAvC5xeJb8b3seB16Qd8GN6HuTM/LlF0j6ZQS5ABRkck2szjO7WF
Ar3TiiE4fO9UQuclZtY7q7Y6u7QYQcvnWxyo4PyjeA51RSBidthIwW33xD44xjSaUNJKar4aNFlA
pM5bnIU5aPBsKUsA7S+hgvdmsbpnSmWY8nqaQOwVUzwkI+pkcofmgj3wuIEns5DQM3Bgudc5MvAP
27UYwuCbi2SAQ+3c3NbRt81NJx2hDjcZqRqBWNfdkoc8aaMGuomXYKV9k8l4tX8i0IwOwk+kdVM+
y27JyBg/gFOZZLCSqp2AeNp9WXfXCGh5IcReDh5liWiaA/3BzySuJSTzAOoVoRjiMRHBD5JuOfSV
yQI1UqcR9Zwh5aQ5TJy9QTU7Xw8qnSdsSooI09HSPUUyLKNfNTV9W8Y9xFf8NTyypRefoxxeNeCy
O1m239+4qrULmB8hKqJjxmXcFoxUGtyEIvfWKQU5z73QeCiKNwLkCNe7iixe5FhnbaHHxk6lmjJu
SBkw92xKl5Km2aZ/uCMOLjYoIDB+xkGl2q+CrmqkqqnE9NbZPnZf/MFDwouiGU0wYBu6ABMUCGP+
iSPN8uaUBtj3yDCOjO0entfSI/ck+UNwViFv0DYBrsAacSQgieAyU83JH3S6Hs9KrZXoqguqMUVG
p1jFyMyzhVCbQ7Jgx6w+r7YwLKLd0wCj2fAFfo+PSUonbwitcckDcsS0JGWUoA6NI4B+ryJTVuRv
2hLu18EPjkL5GNQ2D9+8tsqrErhbK/WU6XlAbplYBU6rYfgg1vmLsJBnx0vEypNrZhf1L3JJbPck
ZAX7bHjw9mLQpuA71Vsh5T9A6fS7fuG2rtQSxBpus+/QtvRG/3pD8X+JCLD/CJTuG7f1/5gNq1hg
mdXk/16JojatRipcQ5WpXwsG0BqYjMXhB9yHpHs+wYlxoinJu8nI9FxHgg3HLC5Twhg0pA7rkyrE
w6mVlGip//AhhrOWQ6DRFhOIyFVrrj8mcA0Dcvs+37M2tR3WHMC2da4radk5zhYgxc6E+c71D8B1
095rmixgvlNL7Yu6mG/rBjybqT8jDB8fojBP9zjRfZ+U0Fz2002RtlrOzrLSeAy8Tcq71rDDWmZA
hs5nXSkCD+A0nfWk3+/Gd0HPBTVjoqrb2Bs+XroE8gq2GHDyMiTnWXFfdRb+oXAAHAkQpAJXCg2/
5oxLA5rmGeFbYBGTpj1/xioBkNzhXgQY1pkWGaX3rWY6N1LOief+ddwvsHuPRynn1mgd5d6QXQje
vNwCzGv21EPmhWrq2MZ6hDuBb8bhvMBSzTHVWJdPiObyMEunhntArYcmUMVxzG8kr5L9BIxK0pL9
oE0JPdRbvwe2qhWJxxiFBGmxXqk6Qvi/xh1WiplmrdJWv+RJ8wlPLdf9YRsqxz+hNyf2WYwvgouF
5iUakRzqnqfz1m6oE69SsEVpkdYH2AgG+juh3SpvN9FHG9HXLT0ySq1ILcdVFC9/Ak6+iBs/wx3/
pfFOBStUfoVyvTFdsVE5E4MeOX6spbF9/lsFNFhjYSjAFU8kLynjZhO5E0UwGDL04rS4jgCXvwfW
Cr9qTbUlSHcFNeGZXYZN7RIQnK9wcI4ZO+ISl+gHEQf7EPD0foY4F7vR5afEEFRgeYdY6WPN9Eqs
1MjNQfE3tpMO7I7crSuHPDc7l9AXX8rHuDxABUQHfyDWUOao0WHiXaPo8QUw9+uiSxRdxOVaRrTj
DRmHD8Nl5mn6djNur0csvmeQytBmmEXbQHGiv/1JpQwEMWBGgsW4HI5HN+3Bf3vAM6w5Vg6cK0JM
AcC2ZGpCwG8iQK3VUaxtOaOfcWlbg6ny8HMz5R0yhZOLgBb4f41qDqkjGY2i3CYy7Bo5OheEVfbJ
zCAEs1eUFLb5xRxqnkREUb8LNjuObpqpHWvQMDHpCu5/wDcbbZaHtTLD2URpEV2eak3+lIXO0Xlc
MeuDgun2HmuiEWER2OkaIdspABctOuFdMAJ6AmQ0h80cLGRuLieY6dmWKLeCYjFMH8ssDofxOaVP
PM8+omWMsBmU3MAjXPnbCR94hNZg4p4ykw+O1KpnkbIwM5JkCo/CH/8gBUmNY0sjkPkWOiK+Om9g
hhYDE2WsnRx4VkfDbzqHUfRsgTwIUFQtfH07YwKn0V1KiLh2h+13ckCTv+bA/oW0Jbyd3qWrSfc+
ky42Er/NadWqEGU5NC24z1FlCmok1CszCF13uAW/9sSDZxoSykjITlg6Vkz/Ro5gz9BYFhA2tAk5
kEmtas9uTFnBGAY84Z09Bzvq2EC1WGs1AiBuFlgKngz4tZCadDjI6P7qH0KSixPFCcxg+3f5mkUl
Oi9p6sYBFYFQQzjZ9S+J1jHRYwcA13vOt4Rb6VwHsk9WbgWxY8Ny3AQjl0D1ubEGzq2SXDT7D5QB
NhXIKCRl0Ej6KietoYQpNLfL2V5r2vg1bn4+aQBsqdJjVG44bYFS9qcsbs5bq3OZ6CmthggXDtpT
nrDiOebwSXjg+VwBxzX78E55QtWQqrX/ehLxFePGX4dAZVsFQLVigdmsa/bxy4zUn2xwtxWRlau3
ZpL8Akht6zw5zdbe8a72jZykS4RcW4DKOK8DGRJFVqVg8FIktFrGNh28dBlmFtkRqQB/QhtFbNqZ
9g+HkH9Qr0nsVg/GLM5xC73olHY/wpQTeNmylEQFhWJv/ygGIi8HCjXuxTAX5UhCyxRuOFKX3lJs
S0UH9YK1L5eCuhnsm87cP9Ph/bOuBUumYqJK+X6QAxUJwIU7gdY4izqOETVJaYJiYcvD7Ia24bCw
E+wGsLgquEdPwJcHO7HlSZkXLCBdjetTJc8HN3ofycd/r9Z7AopWBq0qhO+Nn2Scjeg2e8ZDqC6w
BE4XX3Lyg/m0H47qYErHdW4T/Xk+TFmB4LnbkSBKxydNzVIK5lriFmgg4Xw76kyKs6WVw2NIjSOF
zKFDZvuV2xKqDrXrwx2c217YdANwunpCc1lna87Kjx5D/ZgJ7wMKqrvv8zi2UxH8WTWONPGylAs6
5HGEykeNL32J9GeVhlOVwTpMqKJiHM+bzJ2Thh95UcY3dKLmqbRuCv/icnYkVYQGU0uK9UbCDehu
qtzGuqGs7GAFSbyo4g+qXprNxf6WW3HCj1oSZZkQQrQTH/hO759sctNWUtxQoaoBNEdrmNpu6eaV
4l1Ob3jQbu46pXW4y1TP3hOttmBzTWfF85EYHOczDlIrdPTRc/rT1TJL8KUgiEYyZiOO4vLkK6JK
Aiynx6YnqEa1XNXF0LVaBemS1HiGE4bZ5xeYZdOHyLuEy5DbpQZh5vjBJ4c0FJ6m/VYEidthBh5f
8uFAy+rA/T5nj+8e530sKVS4qPRDc7ZSTj5V+xGzJaplSy4pwL7Pxh0QOoqjawaqpvA9hyGuuQrX
x79a3P/Q4p4SqVWw9zO4Q0r5uFw/IVeX2y81UkLiPudrQ7d/9/cI9IP6pVkhLp2lnUH3cWYBeqPh
4BY9FHZeJ6bo63sHbB8LCmryTrs7c1dfvvwINtwOzjsdJx5urtjzxLfvWS6fT96xj4xPu2F2AVr2
Afhu2GNeYsMFqk4j757BrO2+K7XBJhAdOy4V7f2yEsspH9rWBjeURWJxSq7NQhLOGM71oWFhE96q
YGV+aZuuDdLJ4nNGyJz3gAfL3ZxovIXn2pK+ln8dQWzj0Wqd7iXHZEMl+Qjy6rJ7o69ov2EanFPc
90meJTqQ+IVUfSkuBcjs/8vS0ZnCjxB5GJC9pv2R2W1vNvb2ViUCTilUokwdT/q0IvyX2ylKmKHP
Zua884KbBwGs6xaLIYzzMFMCWST24U+faewOMfvHxL2VwJ1YyOjOEysWJqrF9RQLDA0xv7KnZTjv
hNBJl167RDS0GoWsmP18ii+yAd2s+WXc5+7VrQsmfX4aJzXJNw0+zTQCr5jfNKKK10uo57XQ7VIE
bQJusiw/zmpo4JnGs02m9yLIYwaoGJmMuWn7UI1fAYZ/m0vI3l892xXp30LW66yHwYiNgjzER8jo
Oud3eCQDhCHLRnL82B7RdsE3y2e/yav4/lqn4SXm6rVy5qvImjVPBbrYoUIILLyjLgh5uQn5MmN9
kESkpi3h0GB6yJPHp9JjEEsFXuTH2Uc0lKbm74j6h/mPMcM9p0ZgSxkJijw4pOLf8i3x3aeTE1a6
eyrSssiztrquUTlcxAR5r877Js23k6tpJb+nHE0mJfOueppBlsPJzK6OIG/tWQehh4hHIQFzpM0i
9mmYLKWx/KNWG8unnqEJFzh35mL0o0qDyPnWBXgLd+5jO5mLn0tPCd8RUcjbu+Yc8s7C1jup+l8F
oOCuE56kOS3Dcupph6B3ucY3jBG+ReCWcXmwxR1h2H5bZSRCukqNFFCDiV3GeOPUO5PsXJp08gke
78OoUu40W71OLXbIW6vheV/evAKeDsHBp/v8NSeGgCOd/tQqscZ51jqzBb5VfvGE2aCDzOdJUnVj
m3Xoq0v1TLGKiXc02v/V+rT35MbjH/70voIURzQe4bJ/DoqBVVS8bJSUxtiJrxCadj74EqA2SlOk
n6pmmKnM/hzOfKvck1ATFVbHF5fJoQdv76agNopB7g2D1cH3xQzYvI03Md8uMtl36uQE8BzZ8bb+
CeU4+nogdeORzmjDh1+ecmKyxciw3unKhDY7lZL6UAZMHfBVNVC+B89I+A7j7RwUTh+Tpirak/ii
MBuLLsesJ2NU6Xfz+jn/npq44yDiW0b/00IHVNnWWUyT9bkBZQevSoFJSZHCJPYfxxVjrJdSBdU3
FblutYzPZcJnwJIojCeTbrEqWSc72oxn0Gal0MFh8LOIljdOQkCjTjMSJbzL5yipCIcQjuDvTYKI
yynjdd92+Lmi/VmqRbWloHNu9oxnUIhzlz3Ye5wa7mQ6Icld+SZyC+phwsurmiBukcdmEMxjf1fk
4tzpdCo7c2/PJpGmwOImcnFENXnFcss1UOgOacy3F9/ZLihd4N8d3VLx3BTJhy9/jGs6EA2roY64
q115F66qMI6fs9OP8mvav/84lyj2ni1I8gargNgFUkjtBgu2SYjpwQw7Mththhkl5HOlOFzNOyt+
nynd9hlaCjy6Scq3HEg9I8MNWFDHOwAp2aXdhht8UxWsXLJp2JRGjTHAQwgQ4GrFb3SSB0C0W7yv
QMwHjTEDUFmvY+YqRCQZE7jLT1HrZzhxs5C7Hb8l9vf5/5VBUWmhdB0qnYKQTMG7Z/W1588Bb/Gb
wMa+2h4RjUaTGvp4f2XbO5kVwY4drNwwUs2Lj4+H1QyECb/NpmxaW9EqAVz0rA9wvxqczMFNNiXu
kryCTfSdiKV1IK7+yW2KNXZu2dGOymBgRn+EBKrtBHHS7LJbaUryTTqxfmjxwx4tjWDgMVMWYdqh
AM16/osyUU6s50YOoyHQS48KlOXokfKPAXtqu6SnOJqn+RLcLCP3PViPq5EN0JdzEicfFux1SFgX
iD+gmVk6iBPYdNQdw9S5tdCYOmoRcdMlQA0Xf3V6RQGslONhNxfcpXpQsw5nnorEsCGKAs+SwiZ4
7KCVqmidRZb58KDXBpzzQqZVuFK7/Ker9BoM545W0R/sKUaEt/gcK7Fl8KGCXg+FWOl53G52udL1
cbFLDOztV+ugxMMX/qSyRY+j906tQA9GNdJgXyhvOwxqXDAiQsffqko+HDzO21aBd3xiAEeew8oa
fBKBpvCSqh0jqdv8NlW2UJUKUOE6ZrBlOVpNWFAtMUXIYmNDgF/T0hJmq+ISnR/xsbuSyd25DGp6
PL3D3Lxzp7uRrzfaA+060Kwf6LRfFdTVFYXrSXlyw69wcYuOKTK9aVr9ED9mLWN+NTnmEN8Qa+4B
LPXUI9aFYbJ4uRLtSxeoS59R9UMbBSwqMOuXtls2APxIW05jeQHwzLaMYot4eUVz1FoPLhKzxefc
+nZGbDRH66bNowBjl6mLc5pYcdk70+3mcHLVQwdQVRmeaFbMLWlOQwq96CWH5bsUCqFzgDNYog9c
+LRGz0Ya4kjb4vj9K516R6WPLPp7bJNVw8Ht8+qMzjUNcRbCo1bs+Q+tmxPg7iOkvbt19V852ZQx
LDSmLuEFgStU/eKdm7WAb68MTJoSCOBwxraTOKSp1xeryUNYVX2/IlvXDuFEUuV6eBEmw+1edpk4
eTpSHDfXpXvws/KGLfvnWA53JQ3wuPB4yDrBNYjMSLD+qArdSE6/jpiX9XHzvsoOmUA0NS6lF91i
QJqEPSFJTMLkXUQP9YEndjC8Rgk9bBZ7v25fuL7cz4+qqsY3SYxuTcR9GrL95A+HwQiLTcQNt3Ht
NGRi7B/vO167/iILCkD3YK044tatu+3XxniXe2yPoDefYUBkAR6YK4JdMsFfHwoRKu7eOClNw76J
mNrX/jfPbSr4sbmAUzTceZQy1BnrHH1ewWQrUfw2MI82SFYZaITlEh0mdHd1X+skFWLXyKXzDl/h
zoKwo5zoZu3noahp0Vbtx6Gm2DbiAbOGHSyH56F7P3gzRg8LNT/vYvK4NzpFHIofVoyT8xwOknmM
Ovl7ZOENyIOM2BNYrC6asH6UtFkW+cpKE1oMEe/0iFNWc6m8q+NpfO4vo5i4TCzslEzYGp7U9JC1
76LPHdh33VMdzQIY+MBsn/KgsPY1M5IX6pkgcokEWtSLH4rnKti1D8V9mpeBYY42/GVhh7DxcQWH
Ddcqm2UWgW1fbZw8ziPlnJaONPcXNac+kCV2fdpDua7UV5G7tkzJjMbOBClvFs9u7RF4iWybhAR1
ASy0XFJdjLoOZoo+wT/bHDG94oCLzuMFfkRtDK+6FGGJ47kXHm/vLjn96+CnCAg2Z9inES/XpdF4
WCPNY/Blc56wMNZZjGCKZrvCgXhMIjRP44YcFGwNqv8oqZy9QPdoEtNhRmhv2p1W6J1Ra3Mc5wRN
UP6h0CkpY37y9Brw7O7iHUZcD9ERd1VhUyOloP37J7oXumovRyGadhYDkOh1l93wStqIBe6eTL5l
Q3U3Wg8DWE62eQ4Y4xayjmDgHHopTJnyTJ4yBthxrEwOLoNEj2j27cwmPwqrI+InAF3G2x9gVDBl
rJBP8tD9C3L9gtCp5J/uyrvC0yCcbimjh4igaO9xVMvrKiCZZf4ZF55PJlQ3LiCBj8jtoEjlEOHl
tN/6/1E9lHiRTE/MVMHybMh/FLMtTQ6aDrr5seElbb+BlTchkOYBZm0EouoG5IJOj9UBSNKeyPof
9gBgmmvMniaLtdp/UNlTiPh0d/dXozqVZ12Sorl80NWnOZsTBPwM/fPq/OYvRqvvUOqwK0h9xBgk
MCpnhT2mUmasxTguzFXGg+8RKyYtqLZxGLAXK1e89vS5a9GZbSSua8krW5R7zJ6sTPWR75xaKAvm
+RU/zkHiCKO+zpCgaPYm4vu75/bMSijSZqQS7k2rMZtemMH5VolOZMvXzYCs/YuSQHXDxWDlVl4W
C7RWc1ksr3JygqXMXURqOQlz+WmcZShbdvMQpbcS9J3PjAhafQpiGlWOJIva5Ny0QYi7/tYELAIG
orW3rlFe7JnjJWM+FULntNMuE+hrWqC7jCR4mfNGzZnMEWnUXUxOgq/BJYaw9CUAL9d7I0mNBa+/
OQkcvHjnfbmm/yaGVuKqAlVrZ0b8zw0wAPH/6QdGluUsiv/VT1UZ1LhX23Uavk44HDuzHErcSDyM
V5PT63Dkp15xmJ5o3zGkdf3FdR7N6bDZYXLEL++XnV6T/rJeZjkCqgZfkr9kFWuvRXibJZkUjpMX
lJ3GAYinn9JzJot372odKLkC3QXgGntqZQAiUDdMdLkFbt8SuWtZtqtBOzJxNdzHttlcheMaLg4K
m+bSciTxyjs1MYW4ZLqH07LqSK1i35HZzzZb0AaaNW7K5UmwkQVM+6i9yFRBtPYyVGAYiNYySTx9
XI2m69SEuI4vwbngULUsyqL4RWMUvu1sSHmjcFQeCvQNcGemJPZyeKwrjQczTzawwFuWM1eaUmWi
ofK+OGR1RnaXFs7WSahourO/+dvK3hp7oLiURZK9iOYT+783W/rNnyZLMKmYe8HL9WL2h8ZQihzb
+qTHEdbpgruDbFqWeB7mH7T4k/MPiuHT/iHv0f2vfyeSI6SGDjfU8tFO07JC0qQKMz09U9awL4JW
pZT4BkcU8y914hxUhNCyhne4eN0yTV0k9CCB8H7GnFkHj4jwNapwOgIzO8deYGCKmTNECpuBNAqP
E9rdaJw5XTCwMiPq02S8+7Fwjvxv5Qn7xl5q0WrILRHc8hNbqsE/rM6OiOzP1krQE/8uquSy/jtt
EysdQikD1lyAIMfrp0M+jAuAoxZ7IhbXrR3g9ewIGrKU9zsOhyzaPCxsgxVMiRmfyp3FYqgHwxFx
HvorxNgQ7d3AReuE1I1q6ip5zDR1CnkpjYZmjwkRbvzeot93gndpWAoC6WmtsDYc8YOHDfAeG+1v
uZQR43WeBIaEznD1AUo59z2TtgVrMFDyaQIwGjj1f0tQj9AMnRZnpbmTaCzV5IZFAtrbFQvxEQko
GcA9P3XuZo5Tv//fDMmwmhDCzvFa3qSmHJGefvi+/BppCYRuq8ee0uKM7vqpyrEop9YuBPWK+n/M
tkRDHtmty+lj+2JK3POlMhEeg6xTX+/vq6OXgKXwThNzL+BxKqZC8rSN5AZu2b1dSJcm69FRnE99
H7UjRajlhay19Zxvjo9O6GbAhBsCG6xw+QTT8rZmUMPeGNkzTiKICsVK1YpNpt5Zc57oObQa+R2J
dgxoOoPWR1jA6W89fj31zSoEDZ6KSKK4In7tG1SyrFnZFXH17Z9TxbFe8Jl16dQzTEb+1+dAUdhz
B3HLw0GTr5EZ3L/owwVJtiBAO71RwJQ/vKSavVrHfiHmbwq6ZpolVdQce5u/WdWKHp8jjLLVkGVr
fg4E7ClmsOfe/azVWh/JJvFrUOrpfh4wrHsj9pE32trM2fnFYRGYiFUXgNIbmzpQjXREdM/vq7VH
tgX7VNKRUeAE3gk6jHm5hdituaGay8BniLw7UGie8eyc8aIyrW8R8inJqqeqVoChkft0CFPq16qN
7E7NwJywx6oIGaGj/IK4IlBZb5nm5Mw3+ynEidPWiXgaRxm3+h+bVeaPjXFQIj1erzgtMuYaIa9h
jIxxeeMOr5xWBupbCAUjyV5LPIUeEjIOhjt06KewS0P/HbdQKdB69EbeT5FNLjZr8xFOqhHyqiXH
+fS19F/HbMuypla1ddBuEXYoZQIIrwJcCNqzG8egxAjbXCR/6rTasUNz95JVpHgYPEqhf0jFo/Vs
RMm9JwWjmy6Rc+ub/kt3jqmqOjaTbLoxmxVDh2ws6V4g/n5w3AHuVH17rzZ6BqysgVEV+ebRO1QC
Bwds7hqXU22QUNxlXLoKtlfWSBkJzZ4F+2VhIT1gd76q82lwUM8DqimIA4XzexWSKP4FRPkaJPMw
rw/W5yxNlGLw9z7zX0rXHUF27qPSX//bfKKgfvWXKRwGfC2AHChAYa+yLLVv7VuHuBaVhCYpL0Rh
j52N7bI4YI3TMUfOI1az5fDccpO0DSaMO/AoDsEq8+i6DqqEgnjgGDUXHlGpgKKRdxYLHeA2hjhj
h1Hg8d62Dpu+fJnfs+LbX8sznWtV19hkRUp+VSntuPXbzklFySg9w5j3gjbxDBGaw3TiYDknzBPQ
2JtK1VCxZ2DWuDJ645I25mPREcPr+ZP2UZeMxPBTSYM2rqxj5pJbdluNhB2r6piRt9Dm9nKuMTAC
YrieSWuPW/1jkuEL18mgqat3TmF53lyflUsVbFA83zuHnRLehXhNJjkgClnixvonFF4rJbyVRXNi
BdUArZ6XJCp4qpjTmp12+9Oxej1CNe79AiztRlajXhswspNfbhZT4JkxOHUIPFm8CSlpcDVLAe8i
zypfe5ff7mTytHSSS8DMSb1QidGC6LeTH9SY7WAljWLrmLDu127GiPmPcELln6CgXKat95XDolq0
YXLFP/dm24ZJl4UiU/u3DVrtwNuQiSmUjAtGdjVGlnFt7TC0hi7HJiStG7eh9iwD0xYZEsVN1RF7
oBduJyEActKASU9Qowmyr2kCOXMCEIuMgD/5dUNEkJa0RwxMzYC2HAR4jq9BGTVHyLuKiVjvqVy/
hmgQlX0haT4mQbCX3HPrs8xsb4LbPQFPFrKWBl39bib2l8ss9CW8IgQ7KyaqqdYiaDGaNinfIVTH
76ewc26+k1kGFbZwzc04jgFDlQMycnpMEAvkEDVaowm12+X7hoaIGZBsw8VJXCNlqhDUo55/nxaq
xES8UHdasP1uORDpOM8gOCN5oBJU4gvZtXowqfC/7UMXKvv3x6EG1GsZ0wbBvzBtOCmEczEjYEEP
vq9TmNEzpUtUeTfXjKx7lw8wB8Foxx7sELNIEigCrpkWNFID+2bldqjvlE5B5yjEz4xEft3Sw2FY
XIkP+gmPwtkL9tB/j1HJ2Ov1vNaQARUOpikmDMwlVtZmSA/zCgK/WNDEpwV0/aMM53Q3CTdKPfOL
P9JAoffLsqfZaewLhnVv9HQYuvRb67RClWwFyJAV6JJOdGQQbqpRkRLlxrbKfCvgO0j0QlZvQXcd
SLWvt0DyuZW1weKFcLL0mJU2V4UnfXkd8atAAFDoGS9e4jKcqFZDOND6fv+7rSvVpvnYHdkg805J
ViIRl0nbKnO59DG/PvPa7TaBNBdpRS8HRlmVAgplPeIGsHQWk2osdF+9CDlgYHtNWUxLgIG1F2by
KlEwQWVzn0u9GR1Nhqzfg9mwrE3fnOEauoIDxMDQAZ/WfFl1b66ue0VJb+Cfk3hu6lOK+hud7SMA
NgwDxWRHbPv1vhk3EXCrAG7e6dcAnAe2asP2ju2tw4ysBYFMdD0mz/8Q+etjVMS8vCOfP1tGt166
bujc0WI+1qXYeY46VqBnteQ0ariS7dV/78qy3DhQqd2y65JF2rEYfzE4ZGm0wHXO7KVWIaLwZOky
I/qrgncEDCO3XnhsBf7c1h/eHmJaO7SVBr6ql4AI94yqjLiQuTH9+82jiz3HALGROdL3JhLpTQez
aNSje1fqzViB1GmOOKttU7ePOkKyZQe7D6oW5ryFoB6okUPvdgirFud3j1y/+oyJf4ybbc3K8K+F
NxvdVJho3PofPVSHWf4DMbJOdOqWcxT3rhR4kmAIUMlaczBGG1HxEFRXtRZmY2poe7yQviif6iV4
OL87FuCVw3wFWk2py586T0r7E2Sviify5Xwlo3AThklZEV8vQ4HNFRV3bfoP7QOeO+Y8D8EeyN0q
zQKeoEeVk7/cA2g2Epi04dphkIMYUW16xNP6oBrvhI9EW4DqNzoqnrh8qvkt3h/HY0JPVW9sYerd
FOjm2CEciEfI6XzXTQcOYPrXWGj7aAbNqLbgA5SJgWcUhf60F0djLUpz+dbTZFxG1za8bUWRg9bL
LQa5BS6pLacgWnwTQhGn3xYSKBQLlKFmGfpDNX/c/oSWXhrCnufEB+ZWNIuVfiYKgO8ItGKu3zKw
92D29JvwmVWg9JnXk9eAzWCctq9yEzcSyog7ooKnWSSRtNqPzHvQ7n6JCjnN96h2gdgbzFa41nkz
0GJ2N+1Ps/wF3dkKxJ/ucTICfBZfUJTFFDVLZFAMQ5uqirM8cAzrkvQiAd0l13BQSXTqg4dmt9sY
k8tkVEGeebjgAkG34P5PE8TY46l3/Z6QaGOiZBNfzFFJC9gVt796VoFvtm+BxWvF8J0kacVMwhj0
zcM+lnC73yPIjkAoeuR7620gPOkHx8D2gzmQS3pVYFToaHY5uGU7wz1G6Bm+B1Mqw+qSEhA7bu5x
lRMv6kuzet5GctG53Xk/I34KuyKg0CGu+SOwjUkoV+YzYJUAm2eGEMoQjENWVNu5jijiZ+CxCby3
auG8gWfJkBwhGE5eTm2YqtHTSIrcK2dFdrdaJ0w7KPuUfNskYKpG+oxezPTkWhYkaozk341n0QEZ
cgNi88lF+gGZZqUrpypJVNpXKXx6LbY+YpZjJghTJHMkVC5mbvl4/aGVl2+TuvRJ7cT2tbenHtG4
IVN00FErosCLWOBBYiN2hO1q+h4xsf1XNP5I6zm1LpEJkOdTXLr7Wfoz/SnbIH2b5yqvO7eeAUNA
KoYD1kVC4+o97O2kNqKpNHLsRYeywnfy0cZ6ofOqfdgGqOfhJ5VNKSLjFUGvnIx6zRs5WOLDWi4x
2O9cXZzX2X9RP9NsUQ00OFvL1DYdnSy4gk+qVeKhGAATyXKuZ+VSOkzDxCmZfLc559cL6mM9VSLD
He70YoDCmbIDN3hZgc3zFMKu1cjie/v212PvC1YdEbnpwlHWsY22/vybeeJp4A6lDQ3noq2gwSlE
o7/NSvCzpCataoXXp1a4u4MvG/1vPec61aLu7koY3SXLVJZaVx9KV1rJk82Nd2o5iAZAvH6AAhyB
DQKzeZytmx8P4RRnI4xwBtaolsp/n3RF8TK1BybKFEw6TrPxMOhtGdTWhl4xii4NQmGiH1ajNbw7
G9DjNR5G/p2eCYQtlo5GNiN42tN822CUC6bVs06QkV2sIRFkHVDHhu9fy0NRktoqwranyeeOgSlD
FIe2n8F8mXh/+Hnut1htl1oVEt5f1jQ8dO3uWHqsQM5Hl0zjUDm06VicvOCdlS0WxCVp3PprADcP
kq2E0TGycMLIV2lT/tMktccI+F0T+68aTGR7dNXWacK9iOrAsNPuJ+izRWbWKyYr/uX0SGHx/0s6
bJrSMQ9KwOkKKAhqkhP9ajoyZqv0m3LAqIfZtVyjmHfnAdpNL1ErH4VlgR9f++xqLoJUjzOfI3J6
+FFgAjVEuhV9ofyTY74K569AMXSO01Zykvrf5MP/yAh7Er36kEPSywWI0+00nt6i5dYVNkktuupS
2/GT+2yVNbkrPLRYUJXZMVx/ccnfOBBQCYTG6qfDfAGIRw0C7C3L2boHEhEKYgDjE6RoMZmyiZYm
NVXUs74FTJbfVQEWaMKMh9uVHaVUknaAnDtP4kJ0vBxwN4feIJ5pm2OuXtN7/BSYvDOb5xe8SptX
4cfJlUn/o5PbBJPk3Bidq4wqLZ4+y5SxyvRFWRLFJLCn710/+6H3N5wlXPs5HEr/RsAOSQbjnzAB
HjSJZAGWV93EjzKkSTDqeKbmogZiJUM/RnjTr3fPx0G1BVoowxIi4hUgGPZoia8MBJLRLwmlHZkd
JDySrmNG2v4mR/zaBD8li3ryH/C+gVGUsjJVjGFDpXTcgumju95SUBqXFNGvnzhCAeA4vr5WTmvN
bMPs4n9oY/mf96F8+DHan8CD6pBB20iu9lnOfoDZOu0k8NVh569H0o4z0h/45xF4gWNJ018cgiMM
Ae7XK85Y3wVv17HeDXevhssjrqeM6aaHDMUtBnzfJayyHzWxEfjnUkK3+PJQxs2Y3L1YTRoBRAu6
iuHqqnym+IbSRQIh9lx3QuzTgfPXFk8bDPShu5ZBM6RbPUxiCLUyWbh+jMbCi9FmM8RCiseAMxI0
Hb/y52H6svtZTYR8XG77eJl0LZJLNcrOUOkEXV/WLSO9F7e6JZ91KXPZbYztDP8H7CBW3mXTSKLa
31Uhbv50PDtS8GJ/J9skoax4wF4xlrbM3v6p1Eyb7sOjNqVGkTldI8nrWPLo+DlKqPzVG1K4r3O8
Eucngjnv8bUt0HVmc7i/46Gea1EDL7Z80BGDbJgmfj0pQlkII9c0S/qpdvwGSaOhwwSuh23r/r5C
kF0A8JVh6z1nUcASyI2BfChE8QJYTyh/1AjXRGcHGr+DaB+zjd8vPKnVQYylbnfKPLG9AxCfQw7L
jC6cg4DxV+7rowmVqx2+8to5y/pleu/iWhPvJg3gq+B3BxFPGD1w3tt0CGAhUe3ORomzp+da93Zz
gitFFoO46vNWCixncYusueqku8C4l1mScnLR7XEk8rygHcbrfSigTQzxVJR9Gpeam1wAGhUwGht5
fJ6iNHhH3s0I3YWbEUA1qNScbiXqKdg8YZibuDPS6gqG5oee5eGiHVY6WNK35bZJY1nNhN58WEtm
3mlLxo1lFfOsi8qPGVIshl0Pdgm4jvf17E68GCunukW2Z4YzrMOAuFJPVmK3TBCd2tLydHQsM7NA
XdA4EQuqqbyM4/HGVZdEPeiGbN9QwIxx8W9QyYJMezuusVUdnlFjywoo/L561vpWKY1ueLpyQ3/r
hWK1vJAGzgYaS5/NNdnYlcpfWhP7y3ZBY8DBxZyzcKt2/VF2BRL91XG2bY6EOQxQWTVNTsE1vAEr
h2BvgU77LnPA8X6CRkO0ui2AknakzCIXNiL5GWTVdZ379k/xT/LZKFZqjZ05wPy+hL48dGaO1j9Y
u5M17yVOvOMvayHraDB8jbP5tSftMDTmLnstYUNh4dNSQUHp6fwBfEWUQtgL/ITF3mqGW0m/H4GM
D+rXnw90quZtAhs1jE3x1BVGKgX0CO2risTQLKzIPzPOcTsrjRgf/Kw0XFtCRrxjwFn+cFfCllKs
jFXfm4+aNHyH6ZLVADPzb1+qJdzm9T2quyeGEgnaPvIQ0Vh4NxzYg4kEtbMfIkSg1IsopRny/4ed
U5dAvTSIj1PIDPmKhZi4xqbDe+OfB3Yh/dtqLdfohZJde6TZaQpoMWdi71+YQuKb2GeOf1FSfXvU
ChuO9kTKBd2cmQ+gKPv06McEHHmaMXRVP2AvbmI3CaQdwQJtVlSJjwXmzMvltaPp/m49O1bM8iFA
wQTS0dvqbDUpHPCG2fS+PNkTICzKy6804NxhpNuj0CaiwUnM6QfxCHxcfz9IUd+mUkKC+nyITNAp
XPzJ7VVCHCKMlzfD6EHoZIhbzsKmhJQd4jpUqr1v1Sb/NXRlrST7dSibbTPw+sLnsvlvO5zN0TS3
/+3+G9bSeYBJ2ArOxHJqEh5Zs8IuvNj25SFy/UCudG8QPScO+9duOb+pv3Yv9otDbWkS+S/KlH9l
lqnd/YYzyrkaPvkJH6/NBY3J1oLVGo8ySjJfCIpVEEpn2POh5OZuLSr/SWlmhvD/ywsRe7DijPBC
LG/vAJS6VKciTc5uoYMNvK7Y0+eEKGlvjFRmMBlc5Mz7loZdWBQnfzPoRd+ek726exTk2AD1wBEm
Qg2+XDqYCDlmthKwd5iOz/x8nsPLJqRpTHSgMnO0fXk9GrM33j2YHcBWFLhPDvy8EbR6WZjNTH62
rccsFSnGRA40pTLv/5NxZwmsig1zX2DkBHnEYOCOybeCGtP5Q6GV5pBGHujlB31ru1gWT3wKuVi8
0hAy8di0eBcKfbyVclIJXzxTguauUl+h3fFil3nvVipJiCQN5RdYQAcU2gJSPFc8HG4F8Yv6TYIm
veC+1q2xvRamDU/BQhI2IzkxiWKjw56TqvCsX5xlQ1YaobT9V/wrIUTw0oKM7ZTSLC8Oxrypm+xB
ja2CaQQwfyfEJGRXpWqS0wgCaLIBh9PaShQX+NR7Zw7t+FbR/XurtMjjmNtkNm588XMTTpZMlaJI
AaKJe4Ge+YQbN1OrEbdnD8X9h2n1TxfUzT92nQQNyN4DAIKw2wURgy+iYCMAmBfDE+L2JSm3muCC
cMfrruOEf/7Ca2+PkQXlgId66XrMc/jZQPaeu51WrTOtzYz8GDWBJUBUQNP2f1k0vfmB6DtmIZZQ
tuPbyi8FrP8bOnioVKeeJoS7DATQIZGxbun3DHd9570q2gSjuRFz1+OQTVJQn2bkQIGD4PZ/X6Y0
Z5XtiZJiNk7WGbYhc0rQoQjqUEEQjcYPUJCuzt+Gto8JZ12t8rPO4zcmtC0e0b7XnWaFlFbpXzrf
n03IfocJqUelzm6Iy+Fn8vMKtMBoQfMAcyRl6xBgIHvqMv4ZVcoYZhiBIjSvLXb+ZCXGpSNu8f8w
bL5iOa6bIb7UJuGcreyshdg+RYYTgYc03r/wgptrcKjb1GzFFIuLPppKPmPIvWwt58fjvx15q7m+
9I0D2z9pvGPbW4swXd3guW51qxX9W2YysYeWi2/2liSBgYSpcKkbABc3GxJj7JoIk2tuDarohn54
Chq0PchTuUsLEcKRwETqsTUIOOT4Z8sE4Pqe2kPZ/t/6hJp6V2bxfQprmQ/79JRatVhcngf3pdiM
0inMxiatdkwLOqMxTw9LuuMScY1mjKxEe7ZEjuJZTNwv87G3qaulFiEi+nEFCK/aO5mAvs0WjP/7
bevfX1wsh5cgxV7cxTgYA44URiyS8n3WBBfzZlbYvMQM+pBX82OdrC/KyLii/muzSro/iIt2QRDq
L5ScuIZHi/Dc8q/y1IdUPvcFwFqcqzLLKYLfzXxCMMOkToiLSK0AI7J8A1sX6RLYf71BEQlvAcdp
nj5yCl1vElgGGPXH/0CErPGq2FM+Udwu/hwHNGFgvGvNUD0eFU9ZP49KvGjglo7+6YlLgQnrYtPJ
nWBupmmyuVPEb4aoV5xrR1S+oSJp1b9DKOaEw18b0iYfP1nab0U5Z1kyS5F8VK2y0D8ysyzE13vu
lv0nYARzg+iCBvoX8AOv5vuztwBaQBQTqCbt8Vprb8vEgA2/8TDWfjZw2xifaiQj9n8VT4RDy1+R
au2GavOgCSD7EHIZc2ncA8sUGLDFm2PvIjFukIfu0EIxzRc3V+UTp2KJPIZIfGNT6nrnIGg8CtON
9N4v7otuw1kJ6dwQAB+w+ba88s+CwymvhkMd80b7jyIVqY65gjRY+r0ZCxuBDCQ7AQ5hpHf6dSZY
TtgBkw3bH2h27PgULeR8jDraG9Jt7eDQkXP8ksRyRUaAs+w1Lp1NZV+lO8t5sV29SjVWhnutUjcV
Z6DcJ8AP2BXXjVtHqz1GooRYt44cqw3V2d8UkWpp6FS6VHnAXJRmjT7UadOyaWgLpTx6TlN24/K3
vh9Gti6incbmHZw5I8MUiBsSrqNWumZZOxD16D+G1uHIszAISBvy5shXsrW2bQaFoXULiKaLrtQM
R3L1i0t5VeVf+WU5kypacB8bh1nVptoZdGpHdgTEkebXLMaCR7OSojLTD7RkHKy6GqICO0TW8VA4
R/da+rDvi4a+G+IlQbzSM36ibYrxkUe4w+sdTrOTl5XXP4y2VuGBO2jB+Z867zX2FbkypZUkEjmj
QxPt8OWMIAdVxpDNSX6Dj0zc7e4zukUfcc6np6kP1aB5xGcAaUborCMTZLYgMD5jJknygiuQc4va
xm3Q2Z7Nh1I+a4edT/gkIRcxG6WFrV0DuK67rjqk73vEqcfUdRv4js/XA/cgGoOVEdYK+Qopayv+
I1X+pGnGX0Y2tr9bE/5i3F6DKDxsYHwSNlZRhlFTwxyUXXVx8ipjYSoqYz2NOhnX3st0S8MHnWii
6E1+XTdb1IW0gAnnZqoXK/m4bSjTxPiOF63PFeBCgeAvAQG876XS6e3yUbgdsl1VarUce1uiyqt4
b8K8iDWSXU3xLivBKuX5FQ3g7sMVPywAv2ksA6//b2wna84k4ujWLzA0VZJKC3ic5Ja2drJ3SQ9k
jMXOx98hYJ7fLX4U9oaq38IwXkktgAGJrjKrELzJRFWZYhD1WRbONP/Ca1FDI9JXyCCb2TrO8yBl
6aM4IixhudA7AxNIxmqE/cIkhH0Nppk23Vx70i76E86arOkXjLMe1vzIfBLAYUddV9VeHzYWtDWE
6JxlTot4ejp7xYlX0+p1q0aghHm/0Ef0IXJT+x2Mzj26Q5SlWchYp3TpPebSh5nfS1zuNln+xnri
bD+dStnsqxgICcz5yvKKTzuvSQ/qwI3YMrXw/1ur7ZLuXrlJ5Oy2tGnMwGtlEvpfzbfc5llkiW4J
NDUqgpGhmGwm3AI29Q7QQsyR1flePe5tJLXDl26zLI7C0JfpyPY9NWdiVp82FnYRxqHxA+At0EdL
tG392srXBKeKO4R7g8pHd3DUB+7eorJ9BDteUhjnpuV4BwLtK3Tf3sIG4iVc78vw3GM047PkRlFU
3A8pFE1FRxqj4y+XholQ/0V8iXhw6pP6KUj3kJgpOJg1ph2GnbzsLbwX0Xu6FTYbmo2Fm0dVnVOr
q7kyOH9HqNwE8GVJbg+P068S2aQlfAcJ3Ly388NXFBfRMRibacEZqu0WGXU/jmQ4o7F1sl9Rn1g5
Uql0qzhmDNMGXqK8jGpATEKVQosLQARdSgehTJzK0ERJ525QmlI/dSiXl3IG0lC0s84m81GLw+zk
+B+TT4YAiPrW141yQ1c35nsqL72sBIkc7rCm/6wmwE5lroOEQarDxYP0mzaSQ+6ZL5BtwgOEv8Xk
9IuAhEzpLiHriq8K7N6XslTu7V3RzRQIoH9FhAeQ5tuVbf0ka9aY1VurXtKXQK/0wdtnphVDGzai
G3Ou07HzTeS9ejjToXBNJ/NggyVdiiVt1qX8XdMrpJiqZ9TioiMuEMo3oP9KE+c/oq+efPoGIABC
pw00auANLz/w1qKbyNXcMUwr+eI1J8P1rmxL11TXi4Xa7xQpAZsELueUEVFtCbcsXg2DMBEMcbjW
Zj/ozgMPIzprk/ZvPBd80rsUEwd4QdV7zANrU0u9GRMk+Y69zdUleo3A/ChJTAcq5DbIxFlLHL+j
naJjL7xOcam3BwbxafVNZ7CnFFERZE9iFL+EyR19LBi6FjSp4cRQLlquWthJLm3tGnPclLW/KPtw
5vz9hRh2KC8jI33H43doGYJTfomXo9+WmEHnFMAQFqlQWT3PKEYpJmz2EBMAFUFExYKw0yA/fFtq
XjNUVvDzM0BB5Ey8AzDJyc8bLr2LZnF+i+pXSQxo8ZgssK0yI/AZuHkDaltdriaBMCQ6IgRei2uo
VOQ9K+lryZ6mUovVgxLRg2Oc6ASprhXQ4Ng8UQGk46ZHyUQwiKTDNlBVAbKYTZBO+jnSdmc25jtc
c8wlNLOHGiLrbpsX7EajIlZoG3SfiGMTypiqbfIEKyQdcrRpvEAc41sfjfqoxrKKSILg87Kcrj5z
iwTa+Ph8Ty4uv+VmUdVWrA4MqJz3xTB32HOMVMF/1JkxvdEY4DCzdLStQxzuZc1MWeirrS6dRdaW
e6lXE11t4BViaIx9KuZx+OhEwAL+aD9O5UpyBgVZRv8MCEHT3nvpeZ3VQsFFmBNwul2ojTMRAiep
3LpJ63jeQIg1MZOY+JdVLl8jz+Zz5x2UILhrYpFwZmiYKqdJazaQJ++kJyT/mykCVOqQ5Dz8n6TH
YDp3gSYCPw1CrQPoGNgyorR9omsKtN6BsF9r2+B4JHtBTfaJfN6lprXhs3Bk5DPzxgrhd1T7Xk6/
LF810gT9Rs3M/H3caC301/Vhcrl+hk5anG5asep2tGn3aJq6JTa1OhjkyUdvihA24Qia3dl1C2Zk
mJQvx0aZDEDdUhkKLHbt9vPAIeuN8u1Txmr+RZ70zHHeMpBwMtYN+jEE/00mAmv9kWNXi0Tcrlk+
t51a5JmOe4tKKcSlsDA+q1nJJmyxnnnhIoW2peIpzTqibUDn7VOVNrcKz29rogmLd362MbeOdK5U
QPrbxkG8Z2ev/r7BD8K+H6BzJ8KLGCRzMbui/V7e3wJQsno8R2ExKo04THI8iTiFw+sT5FsW3n1K
Ao5HxN/m/EJu+WPWPHw5T5K/lwXwmJfSoxeU3jnBoEdkN/CY5Uk68cSW8yixPvQZ6Bc0Km1iDGoG
SCIitBJQDWotHNptyiVcsgRED1z+aM/tUvfGmQtgbSfy3U2edwDjK7qPRfBC54Cr7XZZA+0VF/5f
ezaUNeQ7zdP4VEjynzgXuhUSsucJ/MGlt865PyYqsKjWb3xUb09chvp/UNMW7qTV5HpVLItAZZcP
YHRFy9Wb1QDwO0ortSFYpTC4p77vpv/83aCUOBOvw3eVOMyFY1a0SCCZ32NHJQbNoMdhx9oa1qc3
h7nwpXfO1mFAIbzJbb4W9u0KbtbUwKZy6Wo3v9IxRWAptHsJdmkfSwBhcXJqv892U/61kQ1fSNBl
zfjlFBN9zrd77deChi7B73HPE2TVtZSKPo6l33ZxSNm/Sdixnds9oLcekWwH3yn7A8Da6Q/r2W+u
BE+UZLHxZHWnsyrjzuv/um26Si3SwzB9XeCMOL0Lk+SqQeRi2v2vGuR0+iQRkKHkM6lIk/m0OjpZ
OEFP7KPaZfMQ27+g/SHlH+Rn6Lw1K2f1/wjOXZmUVfdlCW85t11auU1FRm/6ng+qLurNcXW9TKwc
/Tfe238zeBSqyZuNki6JPUIK6mq4RQZwfVkPLCmlqP2RoWXpxV3tmlnG6lwpA3yrm7JrWH/0BTxb
DJt/PxhOYeKdwyr5BNmMqS9PEkRm+I8BtuK1ixX2buOVroD74lG0rrWe3MM/eLAeBiN9WVZth/aC
eWURRUgOsz9fnPifo783OZvzD5Kaf7lts5zdCat4sY1dCPRtQyb5GHjqcc6X7qQFBWaNg3WhgXYz
8xhjRqvSBBjDhNyARUjF2/Y+AD3lTGU5qFgS62I+RgKI9r6tF1PhMXp3B8cUdymqkyLroP7wkLJL
2Gbri+DaSummg9tjelPxmQWCcNKGpTuK4SNl6lwZ4EK2uTSUvfuMITStJwA/Ibq0981GJTULEKeI
5cbgDMvqr1/AYhwONBN21KTp2ifj9qUw+nExyWqpkZPUCEEw6KCvmIm8gymYC0apvQ8JCuDo/wx0
4YqlMctg1vKMzYcPehuKHJ8gczoIibjhQAAdM/5CStnAT5UVwWHFvBJmY5FgUL0dyS3E7OU5Iod7
VIRrewkPgqJPkDFM6z7AWZKWnq0caG+DVM3+ygTJmRUvTg84IkYRglfky7N1PAM+uQV7YXWxIwUm
bhLO+gVfg5/qaHTAxYZA8tsT6QUH5vduiDhifrsSeFZeGjJIFLS7EsEw5f8IK6nUwCQrIyOethjK
Iy/rv+lnBjILmcyKbh+bK2YrYHvO9cM+2Mun/vxB/WXQB/9Z//o6XfBAtgt9nKA/i/7D5l4WgG4y
oFwyBDs4wsiFJOQAuYS4BkTz9Whab2bTIJKPeLjvKbcN49Jb1G3uD5V8N1zMWKubrxbKD3ojmMYl
T7NTiiLqcz/hhd2Wpxp4P5gudsQcdFGf9pMjq4bYP5nYyMi5mHTxpKGBKYY73iPm7TPjeaE0/387
g0uS8UfACYWBjsEFnvr4rZFxik+QAiwmz7puUnvP/W4RXTJIXQqcHaLDV9IKMuopgAy3BwXeYN7V
tSxWtKcLOToTgEgbM9ZsTNwgsjgqnJLiUv5rOsABEonI8KI9v89KtpylOG9zFRiA7fWmjmMbEifS
9W//UcxOGoDmYf621/53w5Sd/BQG1LySF9Amil3dK+1cPOKX7HppE7LK+EUSvSWHFvCVVkizG1Sf
6xIjU9dC2Cg8Z5zIdgx0KX8Kh5D+tlUAIj77qsv/Fbdmof2dJ5c8SHKwpg+FuXqmhNSn3EQnYhvR
RoMGlHXxkpUVe9yuY7cS5rJWQVA6CCHT9v/74eUTuXg0HTFPuWdESugiibgpult2pDUkiq9h5ovw
yQVdPM4Qo5frrlOjlkSfqH+RNnJ0R/O0CiSK5pf6JPhnlgrgygn4dxly0RcWcEd6iFPe/iQ/N/cM
3SLBZwIQLbbjCdkxenkBtAh6TRUHRXcQoLbuMTBIbu4xuVfD1/5FWjxc7SYYPh2WyI9SGLZtYCmM
RiUAJEmj9/VdCMatgUa6obYBhljwbijGPINKHHt96Mn//+sFA5A69o2XXxJN83WbEVmY5gz9D8o4
I+N7jsJv+dbIX9lR+o0nN0fUaBjvNzoNd8Aoy9O8drDeNnKpNuzefF4F8W4uKHiZmQJn2r3NBHMd
9b3JFF8YvQoQAbbdRQEwkuqNa1JNULTbEDyPr4Uu3soa9Paffk9dNtpaytoMgZhx2tcusfsN2A4o
ZfZ2/gmNqPuN9bc1zsw6ewKpimfDablHctdG39Ltnrm19b86eDuXoV/nSSTDKIBA+H0n1ardkf7o
648ZAX2Ew6PDf8B6dWLSYwt/ojTOzGILLCkQBeIxatqlHiuHG0zC8SG7CktQ3oJ0/ec5h8nJJgla
tax5nc5AD6CfTDWaqnk2jOqnOQnjb3wF8QjBOQ03xmBjhBzD7cdm2SNqrjis6w0o7sghL2EO+sdz
dm7eUVw1A97c/UMXyjkiVtfBDU7jc++4f4tJQQpPObx1FlizKz6tGjjrJXiNgR8zxJclpSFsjMZ8
GBTocvgf8yF9AjsjEvqsGkC7dZrZdcoh1mzCRbumCIILAvw+Wy2gTGWwplF7MlR3qRBq7j7D8hJh
pOGeZqFKHCcb5l6eOL7K8uu2WJOqTZ3xxrhxXSuTw2yJw3LqPSzxemvoU/LWkVFjuGKLDEKeBLrj
7CQ+beKc8z2moJ75Z/gRgrup9DVN2P5Wqu0vgBbjskQQ32JXOusk8IDHNPXOVbEIEwZNz8HcnJt4
96dOxbGeNQrMYgVNht4RzrObOOFWBYA8B9yMFRTnZf+CiiuWOWZm4T/WeF68htOC3p4ui6CK/n0/
tDVLNpsAegGWlfvO/2Snou90X2GhLmT4J4RYVTK+06en6oYsdXsk9K48ZpzrTnJnY+q5IIn4Ktox
wMLhFakGvclvHlki4ilYgtVeG32lajpJmk+XyL2IVBYMwI5x6cGby8zwxHxZXUTA0CW4/LO1vgfH
iIoy+0ZEQTqJNh8xy9hmaa/fLBLmFYUJ48N8Fz9dwWDaJC2zqutbGlk9TOsMMDRtZl6OVz1vpvWP
MJ3EyaWeaz94ZXT4z7L1rikXVgnrezjpN5jnoUAFoLbM+MfWKa2hj+cylI6Vtnh2KKXlwDGfvG2o
trS6XMdPlPJZYjQhDzz5omCQ9ZlxIRUk06vwDVoSoUztDp9fhvmyLBzpe5dQQe7Gc0OLFonH+mEf
JYCScgzkAiOW3en/p80HhpmOHjcS1updic10oA+A0An8RbGHIdGhUmZlEjMnsXPTeV6fKyb9uqm8
Re6FRGqYl7qs9lHKumO0qEV47GDDe+jZmdpQtRAeNxUsCsOZYTA+0hG05XLxSl2Y8Tr9ZZvfAgi5
PvX+Z3XFW85tseSBZrrncIHP9Ufl9ITnD0CN4/eg/t0FaA17IAZtXDqnds3YMNnzcXcCpighjBht
T+WpAw/AZduN3adlADJlDBkt1+UwVXzI7E0xvBgFf7ALLoC3WpI4Cc8WQeCxLJ5MTZYlCqlneHqn
EM/ag84zCtIoN2PfhU5PBwRljYbnb3kG3FQcQwe4ElkT80TG3tfn86QrKrXOSFCk8SEh1CuoRemT
oRZNIN+rHV8nvWQJ8g7J2wHp1VuVOr5tF8+WdzyzOhzQdZ8a3+pISgOGhd9lbmZFuYp1GIRW86Y3
5Eu4+DHJb/+sqwAMguPg6tDe3bWSw8Sio9bZr/1wfhuLcpEevP8IgXS1epZeNusgahz96O/Ej9AL
katnpuoyvQAXqT+hTFO7HUUF9Zo5bCDBkU/OW2uFPS41znvrIUcVpzoIRIisoUThgNLP/4vdfaPX
NtruCKATH73hLqTmnqzo+kodvq84zG+/aitj6ySr7bGDs+fZsUaOI2jNazerS/f+g8gB578kD1l0
Gd8Ec9l9xgjEcEYUF//dTzM2TGe8yml1PNN2QBszVIQR0khJ+OpkIIs2NabWLFwPrOhKPtXf2W7i
nob0GdV70mey1pT43CfcL6HNHU5pBNkxyoqI+1ltWLA9iU3FmrSt+DPvZ43w/ReU1yWtq38Y5Uni
njgTpp+iaa6eqzPVJ4wvveStdB/mk24QJ0kgpdONN1tFlRgXnCUFA126wdStSopCqMiVm5myBAZu
eGU5+KaJBM9tCrs4HaYHHtjq1ikt8rgWzq8E3OpYjNPQgoj9RL89ebveivKbQiueKUNPGgX8FhsK
tHP/A29eWwrXigQO1Z2PwYAyn4NU8cA9YjdXwR/1mrgQcPPTu2zfmBXCerEn3k6vZbG7cnFEAEJx
5z+DSakcX5DqccWUqrtW68aQjDN0UOGyp4LYzksKrdDdwWX3K9fyF99JuwZtv93BFBJlqpSblxkr
rdCRPEwUVskpFfqLF+KXX9WKfjhShCz0IUzyNKLhmlv/15vfeXBsW0MT0AEil3oJ2ecQhmVXXZHW
paV/mZFwEPoUtB3+mOM0EfnseRcxF94KaASG+j/7N0ryAS2gBpRpPKQe8RgEZ7BuZC7hMQzwl9m0
Twm1+kaZjrRIq9HU6tTA/AacqT6L4d1S2lQVHyjcqd25sxgEjPaLWOO6GFJmdbFIFxpFSbDWcTlg
HuIetomAMZ4eJ04HG104tNjHpW1iIE943h+zBEiGLd19q8fRwOJOWWjtUOPA7fmjbZ+clDpG/V1n
Bd3h3FlFGHcxvXIClLE2gOQEV4dgcuzlKsFXvEJAZUmsvrtiMY+NWScmRemL6hK3HOM+SStgJzhv
4HTJGgAp/DS6VH3+4sbo9lWyObLAJ/leW1bGkyjyvMYRCUqmhqqMcNmjPwvj802DigSkPX1q/66P
snB9+lvGdvhsdZy7WCw7jTih+0LrCcQlsS/Ry2Y+rHmVx5CTLDfg3cqQS3wsr/xANhMKwPJ209CK
1CuyQzMWNchWhXdsSQ00SSGEtKvIBIriTKMjz/334+7bxEvVnc8dG9uETAawkokt/UDq6Br7lKoG
L3qn9Kwlb3Dgm2ctiC1j4FeP/9aLNhAaAYHXzMSoZggzC0U83dLfD47LgSO+g7SNR0cOP2rIPx5Z
5xA2WLRMiLyFGlBegx3usMLOWmHa+JVeT+F/n9pxMA8VSIbHrxjiF1ApSc9/XsaHs04JvnB+XyfR
LwNadBDRG9BAoTn9pdEXNbzOi5iWjPjsLDSUHinxTQ4E1UbSvVvKL1/dCkl1Y1Ogq6QFUWfo8An5
fpkbM9KidpCfkw4sBgVPussMhaJFqFCwDfADDAqIj84TMzzdfOF6SJ1HkwK8tAoqqUykEMsW5uOp
YN5H9nyzaGE5ookLeDZjsKLNxyNv7hD3InjsHDReFqg0NKeHDBHS+zPYvsg3sjyS9hQ/4nHidDrK
Ux9aUI6HxdOCpEYFw1xSxoFjqbkO/xBMm4kS5nQGlJAJL0kkhPCUzYO05/u8lKmysTYyUIKXugt0
4nNWW5OEh6zMhTaq8b2zNhsVd8utJ+kan7g/HOxbI9JDeEn1dcngXbjM6IhkQ13q8/Ke4DRRtnFt
13irRkBOWyS6YMToXX8TXA20rlKAtMv6DSHfjLAEv8edwhmmK9DzDJlvoYrCZjMuFf8yDZ+AKE3s
4EL3pCEfQvtQzZzTdjsSKOgcGSe22obEB02b6C+sdx6pvOSxesuoxW+o1Ol4GFU3eRTM3G3fAhY/
/oEwHFaeAuY4bd6/qCQWrcHCVKiABxSEqetqZ4//x2HLUyiKtSZFS3jh0mZ6duTay3eYCy76AFcD
WtwOn1xfnyAMM1J9Y/JyLTj4tqn2v19UUIZr8Na4c3FbHuABaX4hc0yCVWH1egpM4G+ImZvYSDQX
LeCZD3EhDqQ8MfjNyrK47ESLsabUEet+peNEA6SctfsltGcit0rCNgIp8sgOncKgZYkpbOJcB02b
KlW24UlrHiuvV3LwCYp9iUBfWMGZm1PJGxMk7/RjUhviTJbuSdUImCms5ocgfGwVhoxtqtSwk5Z2
OQb5xS3+59P87f/chrHYspDBQcJO2NkvqDp9x+CK2bqKyE0ZBZUmi4WLgeI0st4cyw72Ecd6j15l
c+xO9aurcmW8cmzt3cVggXrmX4El/jzcplr8PRUg0Wy4opNZSOllO/XSdxqgNXeMhhFc+JjfcKqQ
JSITG0mqEZAuFvXRe+ONEvxJpWbjaSKpeWjvkGxzXwlNAc/Jc9d8bUAB1kuUKlj6Y8Mxb+9DWr67
TORwJKlV8KMWBZq2qzLEkS4kLc4iBQDKvn204wlKYpWpYSjRVOWTwv610MPe8J3+c3MYLzPYpnX1
mr3LT7nJyAk458kBvcYWNAHlh2iZyT3FAgw6v5RkyMbAF4sbgTHkPRwNodXT+vM2Vvvr9EfmxeqD
gW9kcoqCY3N+S9Irwct6CZb6dBbc4TFlQGI2iUHuynTKhIh6mo9JRyXtvO615AqKKPcz0flpXlQo
fBocPOLSTvGdNyoCO3DvGXCaLDFgJvCkQnMM66NfN/osGKBZScijQu5GLgMliNfn0Hel5vDLUwA1
ZKwQrw+N6NJsGTm2MfHcEFDd5tyKox9hmX7q16pO/KmZJwsQ2bHJr9/9eAyeugfo5siqWGDsZCVm
9ofxe0+s0bCtWmw4aGM/kn7+oKQs3CzbIwIjj+LIOg2lKg3RkCzIl1Yk9/hDDhCTwrQpZm/36thP
CYdtXeSyWKqWIdwqHw1yI8j/3CCkkI1CIl8j7Ejq//pc6ZvDIvSyTrlFRP5tfUK6DQI32q1SncNk
bXN5BaYt5VIrJqcnGlYEgZ6t8LHt61YrSjBXEfSH5I9EmrZfsvNIu0VTc/kKMAURz3b++uO9134F
myQM/swwqHqXnVRZ+Gul8lV8j3ZH06uWZe+WApZbFtWTgsETPzmgN+qhVNi6wP+kxW0uOh6rdrDX
U7L/cnKoVEQPbp70g3lq5TrHoBxg30oIZJCgXm9iaUN2GyO0BrzRv+mvCan+c3WUgyMN6tf7VfQD
wfjybJGwijGsramglDdpQR32T92Jx8FUSqnJzQeM3s8U5dfWr+8W5OQrqEAcf11EfErEO2pxNyys
Hu8l0MQ9DZnFQftqKva+MSNq7gQSwEK6OX9UQ+hTqzk80GJd394nwhA2TVnqBoyqu+54sxceCF+f
nMUeA6ZqLqNCMG9b83fxBdL1wZVYrwS+DWfaWb72slIlXf81mbNn7u/SPZRDvvb/vPMGw4yKEctX
w4Pw5tlaqF2Ty6wGHkozOckSifNPKi1TloIRrJnr0DT4whBo8vgQQeTTPLgNHzcfx7zuNxcmGxOQ
7zxSss8owl3zweZkxhvrw98z9tYnc7mJrKOvTPUISXBMoKBfNYZJS2UUYqbY4b/gX9IXoWPfXAHJ
H2btvAEnWjUUaQ0NkqjlnrMyWDAIREWjw926kWDc38jCeZcjT8vdKPFaXmze2Q+gFCSJW+WRPCMz
4KoTxOc+06d9A7GRUp1t3D0GbJHyew4t9MgsVxB78SaDztsN6esp1W7usVYqUZ4+dXAC0lzeD0ZZ
lTDzP3Wi1TVgw54CiPT/4P1nE4gMvl6Wp/dKnt+B8e9xzS/2mimEWhT38i8vL69qFrCSuFIpRsTM
I8HYsKDpwhEtPrpdiDz3kO2wGd7AtDG8rEk9tK+WAF5+2Tj+xMpHKCwEllxZdcATgQqgMFqYosu7
u4+JEIn0n8w7N3S7X9gudqeyggZ42Rmz/rcTkssPVgF/Ie/LBssjLyBCcnZckhCeSJmX+qwnsY1V
YTcKN9MfL+V7t6bRif44AZqEFjVjeiAQsVbKWxPemWBgG+hYwGkDQ5n7G4Oj4lcyMPWR4h59odJd
yxK3pzLHsPOK44DMTxr1Jr21sDx3GGmy5EzuAaK60Pa6o1uTpCsStPSpu1+iLxNnckl06LEbB0eT
6kDiaNBclvSO89f6GOSWO0fQ2fPHJfCRu7o/3Himkw+TK2wfHlIjO4xNELfrbllG/JsYAMxQ9x4k
4G9OhQVv3tvq9wdZvY+GTWyc6HkvKOM29hOquaSQQm8FvDzthntnselRUgYw3xH9Z6dMVvuJt0No
AXi+XX7t+yZ3jZDpPgdMNMJioBqT0keTE6Qt+oC/U5TkCuMbS2GLd3vQxvOAK6C0/4Wb+wpJBp03
xbNT7KA9Yg22lsepuPmGgTyMhmg5fSgOWyzkr3UGOolM4OIQHJsafN3QTw09lYfstEwAnDdlbLKP
Hc2xX5gBDTJFyC6cQg79Eh4/C++4Qk8dqrT/37HBAUGfdTFZIEcMTn6PIjruIiFVs7vibCK00NVY
zCU7Oj0Iz9u1CjD8/DZkI0U/rLRNUFBcVe/22je4YaJGgcGqCq5CsOzcM3Q7gmidk1m/gJjcJ8l9
aGrZGb6msUP5u5z9lnc5CBJCi4wEhXw5O1bqYQflkkbc2oMZBt3lH20NymC0F6YzS+gGJTKZ49/6
r5Q3oyKyTSzaDdgv/eZIwNOBCJ3n8mKDKU3HcHBN4VYbUiCFedAAAg9zs1X6ZBGAS/VwT2nyaRVZ
183eEXGsx53m+3N4YGWXVwmb4tfWhRZv4Nq/Gc5MmL/mTDu5EIL1JK3vPzVet1LR6APD9GdrArwc
+tZsowUsSILfpWSK3yQAB1gn8V1jGNbvOA96btOLi/0sl+EGJ5gcq9b0M1Eo5/8860kXU1vd5coA
ySobd3Mi3ZEOiQmxjgsY9PV+jzuik7bcPDQ8v+1R7HB6skIw5m6Jx8NgXPEZTE4mGLakcYPEC17v
+K52VOMWL1sPPvigzWH0DT88fGKRaxigzszx3sJS4ifrgbzlD0NKajA+mx5SLPxf2Qcw+m3n7CvS
zp5GlqFPCSUERRk1wKR9CW4j6Z8NyaNaje3mVE0yNebMXC1USnTh202rHRtnKEKoMKbqYBsX+T7C
mjpvS9jXb3JatX4miWZjRpTOl6i6z3FaxF+YKklSXOEBUxwUibMdbvtS7oiLfmDanK1xlQs+Ehg6
+ANWl1PhMp/rsLKZz6rB9Hj1NAQvGibp0MooUZ3cBxVJlay4NI1PVnBBhgBRzWTZWNEMcXIWlM61
VpS+irhe3EYbXjg09yEjpR/pZQ0aIzSEzaJqKEumt9pHeY013TlmZ6tqmvFIrcgc9DzauCyF0sFz
0A8wdrIkpUYbC9fB8AVa6290xf659A/663CIIYklthp8RbP50Gsl4/heJN7lonAwFDr4pLpf5j/7
7j+eoaaB3Nh5tM0KHIKTphyZSmynNXIGas8h+gnOWjdSDYykeauPEW0TYUTk4zN5hWOHvl1XZ5Mj
PYO89P5gOD5rsqISm52qL7jU73JVsgRGsYkq8WFqU7eEITq4kjjwM0CqWCGqdthVR16babGnp0A9
H4klAa3IpCEANI5shqIHuUwINm8/mfHdHCIzs2surq1H7IsQe8UdxdiwlaEvf0zL03yQFC0Ck6ji
LQMUfbt4UdP+itE4etSdTw+EnUQMwSe+CaiMowwqsYilCMaDlqprjXhmlksCqwIyfmGi+Vi6HXB2
1PhiCNZDV+JoLTOrsbrXVHqMckudv5UkZU00i0UB2VLSI6vfbxF1bqljeyOOlKqLOLDZ94eHFS78
JR7KKGtCwL3nTfF/+Heg/8ipHqplFknObw/nNDjvAXERcaxBrxsB8k6FLf2mjhXH5BSuoAmsnh+t
UiuS4hXJbMmVkjM9mE/Y1MBasj4xU0UtpPYqFEfqZKBde00+O2fsak1KWdzlzvh5nqudltUA5IqG
6cVsrjs4c1rQMI+l+KpX78CG7kWN62IZ0IMePfm97E8FKGtk6dX85WCDj2LBYDCW8UOdg9hVA0s3
45BWKr6SxXfVvs4QMjJ1q80iHLYWt5i26T1HwRf7bvVYKdrP0E5NH4J27QQc0b1nuDgvURngTK9V
dlLZc3fYTC6Vv4eKpoPstbv3LGgYCGjwHtQAk7q688iV9eyZZdbGLtK3KxDEJniWgyWz9PkBitUS
6I0eVNYgSFiOdZHQCT4WpkeqEmk+BqWKvJ685GedURmD30E8SWa3UrI7lWDmc25St7KnGsTVYinX
jdq4sBqF5GLsXYRAACKN5nSZzmiu/4lcz3bjdxgXQfraNpimCxLcdJ3B4bDyT4Bvq065hJEucloo
vnEKY6/HXLdxzF7r4RH3MPtBO0b3Sh+eyZLhIwm6VWq+vqu7HGaa9YEJd3OTpXfNj+F4hEgIMbA/
Iq+KM0fSt13DbkDx8VFl+jM0/nz5MA/LAHs2vp/2y+vkzDVnn/VKIxDhIoCufzMn7oo3S4EyQEpP
pxGjFTjCScH75sYDQbeUjb4RdxLrwpWq1IyB/ccwg7oE3Y789Jtsl9Q/20GyvWcEszYn2nRkwznU
MclLTPidDW47i3Rw1OKnUEp2J2JqmFUNLBP0LhJK04Da09Xk85/GU4sz8bHpsRcABgv051/IN5Hp
TpqWe61vuXTIvZNMN12NiApTn7QN30QnOFesflPqdw8qO4LbSCscA5qnn7AFab6mM62Gw2F0InKx
q8cAv0Ptc05ZLY4mw4RzUHPR6M48eEmwIrB9zd3E8x9M67Mf57uw32KrN/hMSZ598hb/0AlQrD5p
9XvRiAbdyfhZNm6Gh5zEKDkoiFv4IUg/9M9u+i3jHMTCNyXVTzE/+FvSXN31n+Qa87SIkIIH+CK8
Z+OJOy3mezgmxOih5MAY4AZkWotLE9b3zB1LAmLQRvcJAuYz23K4ax3QJKP/xTHx4yy3dIA5udTY
qKwvxIAMxaihL4lPVMD2GQrijblSnEvp5u5VyAed0TMZShpokKv8i1qwukaRGM4MpZ4imOPHqW8c
K4Jdh/hTeqRLZoIOAdEj9qqeYB3ttVc140aMr/986EMm1Qz6FqRH28PgRMGB40YrXcaqAAi5UYpv
1c73eBrIZNtQBmr9hak1hrDg8zFnnZoyBSBoseiH0DEcPCU5vTv11/RZWhOHtcNXMPlyfnhvgaP0
lDbD+ZoY2vxYnl1p6+mQk8jnuRQEscYpxRabjNe4bbgvic6DkfRyZbOHOPvNSC567SwwaQ5XQL9A
dCIDYC2ZrtwQTNFiqg1ipdeh3bOR0Fc+bNoZ8GSMyENWjSbRvcvRGJw+1QSwjV6kxQABc1yMwoel
KbT/7uoUCtAxciu6p/yKAYUE6KgvTBb0KNiaGQ/1J/qrL6JALY6zswZo1Rmum3uoWmb69dk2/E5Z
lATHqs25JqIw6QVApleFmfwxGEIIzURIAQJA72nvkWXu0KfpgBaEjZJZqfil9uOfa5pQex9Vsqgq
vS83KLSkI/rC2LFIqE8o8Fn1BcJCjl+XXk4BMhkwbGWs/W9V12U7lWk1fu1ZiStTf/Bxybncp2VH
zPI258qLophp5eYzu5UXC0AqNZR48/NSURytbZ2WvYjR7YdScCm5vF/h64iO4AkWa64k+Oe61chu
71rNC4SEyupK4n41anCQ8FVtq+T/FVBTABilBdSXcQKy8wOuMfYnR8OqVevTrfRp5crhgkjZvIIT
N0jxsk/GQEf6+UFbEq6tmdsP4smfPRp7SswLcv9WuUe2fB45WSFiIUEbt7snR28MFG+wF9kcYflg
xQ6pJdn2zYM1XibP88i7R5DKIZ302z2vUgFRwW+gMlsK1y2h1sSSfUaDuWMcVn6BJvwC6KyWXCuJ
Y3pxl6O8ACquW9mKeMsg9U3tQNeCEEewd8C5+EaTBeJMoFRzG1jFhXeJqIttK357/u2SmIuqUw5P
hyq+U259PLqlOey4A0OS4QLtec200BH3AfK32fo452uOz9luAssN41Tf6EBfTnFqD7AjpwQhhRA3
UZl68OhyLEuBaw8E0jneufIJ0WA0G4EYZ0G3vebMa9sU6Xat8cQPKWLZ6gCVE/PWmqQgP6uncx47
eeXj0Wcg7oWJ47/XodEpI45Dau46A4RAO0d0ZKVlHdiqxUojncmSTSt0vFKhcwEeQwfz+PePXOg5
N1q3ERx2IaYG/xWo5dNs+GWm0K2zOa3147Y25dSwb8PNjnT0hDRabOT0oaawkUePIH2UaXDkQUQF
oeO5A7kPNvynNhW6F/SWBoKJP5lY8JyQxnSV6KzpnUP1w62PugRqrnsg+AmIm4fZF9BPSEnTu2OP
bl+4Ev3/LSLUj1JQgfqrHPYRsAfGg5s7dLh81IvDdBlPJKZGDddl4aDn+zE+R4sWbPmtXRiyNgTn
JHXU4mIl7c9C7OdbuQYdYOrqP/33v57tXuV3+4SOfRf7cgBIK8czJAXm+apkFUKqsdEN0z5ScCAp
NXZ7GWAiOSMNKFeGJXx1wkL6XAJvI/K0ej8m9R8JuUhJdX9DZKSzB0i9LldKku9f1DBYi3DJ8N5k
bJv+JeHzauDpMQpE6xFi8WqGacLo2AZSDUe43Dja0kPjTpHKHkbXwVsqDmq2X3pX4gHqu2nHYZNH
HxTMLge0sTnm7tGki+//lglTvoshdMi49KMKSW9bdAur08WfTBFwurblVm7fLpTPfzF1pvV1XIax
cL2IwK3RjL3+ZpQ5MIVMGNSxB51bewJ9Hz02qLs452p/+BGCfQegB2ppqV0SqZetGW+33JO49RdD
feSnZLxjUW3WXKezm7XgQmqRb77TUxGty04q6D0TTOrgpkU8vgS/B5+58Ku9o09N+Iqlkkfk/q8y
3cbpMuQF1RN/HsyGlp0YD0N2mhNCc5g16xViv2e5iTcdMQcy6L0CvigTx8McEZuquDCN+y6pb1NL
YfkhQ4fOoY7jeugwhm/bzXP4pQ0EzYaYaWbNrSCWenJECi9zwUrI8NjDTpvs3azdBjTWisyW3v+F
igNNVW53+0J6c+LjM5nM7e9z61hmkTxiWI9038RZ93iTlGq6lbL3P+aR40jv7Uv9Ep/GtMycEYhO
TbLHurIO5M3P6ZL9fSOv12+CidnBdbVqkWEPuWe2PshNTFHsv3Xkbz/sYe1LFkypVgwe1/zsHwwg
obKEbUzoGSFdj+OD2uN8LwLAeoxXWhLFvHMcbnuqz4pfZo0oQJwWfyAyTFwo0fj5fudQDxGIR+L7
czZhOMXm543SpbyiGA4vWRANwds/AaCpOYwRhexBP8yUz5F21RlQ3xlz6OUr9IxMyfRNM9b3Ikcw
I5h0EC6Vo1Kb/AZlkY30W1191WqMHxk/Ousspk5FUFX0n0s5gUbeH9ANtnx0GvawKWri+h2XIoRm
YAiY0KwzPEaDsfHdA3R8ijHKLpyEC51SDojsvbge7yS+Cdt117GAFP5RN8ahkEWDQbZMli8hIEhR
X6/tJwS6u10x0P/st8l11471U+N+WsA9TUMcPfnJJ9AJWdPjGmA6PsbLeEeMOzst4x5HV6D5CYSL
yZklZCySX/PyQUQxyNA+HtfbcpC4d3u6LkGrBD0JTQ41Fa6c5ylwLGCuTfJFFcz/dgM6d5y17g3e
Nz669KMXn0bHYWa076xyKEIzpLDRmpFKdjyXltyX9ycOQIwXvE4T3oxOi7kWez/57vU3Lyz2S2Np
T1DFypKDRJZcmCJrQNtT4rpDmMaEXVwqyOSvz3NSUa225rvkKgyMpNerGjzcKXcX2MYt1/TpkAhz
DFwKDHXaCLzPre6m8T5Zwzy4t3Ur0iZK7b0Ii9T3cknA5Ba2bjc8tr717iqmeBm2ygUzmrxWOPO0
IpyGMyrLlcZL0DBH5I5wapcaBtMX6J+I9z74ridskM9puNlGbgf7Ik8CO6njP7GlLB+ip/YbDu4j
9uHsvbIeYqfftIHUbN+/MicGJes7GYnTGk2AaaQc6eHRvOboTiZ1eVpcvbSe0/+ngOq5oLttquWz
BhYKAPWTxn4CZa0jeNAhIfoW1ehI72vys6Our3uOiZiAOWh/LnL3SmqmemuX7e8H9sppk8Du7Vzd
J5P6Vkw5Jx/W6ro8MMEhwbKSqIbhwM/w/7ZKpy2BZZ6hewhmym0iQ5OuuK/3fbDvf2cIb7RU+BHX
lJdToaD1HhQIqedpudez28afUlllA7+JZHKqzvxZ7Izxy4Ce0IgaGzEL2Sq/M5l+Irvlbm4kRsdp
uJgsqFNgPXQJHgRigLjO3EFC79gN5Z0km88WY145sNs3O/YvhCQSvaqXvtJXNzmxyM91iPnVvmP/
BLfqYYb4Psuh1EDYI7qTcwpntx6qN6yaE9ZPa3Co8mH+1/a2JCqn/SMkdK2QaWP8KbPx31Ii+hth
Of9kFDjEuJrhJgoCIY37vLXPHhR0WWLoCvCzGp2I/aAogYVldsDGGcaV0u/1iByjCCAVL2xwhPMa
VWMUbM7LrsLGfBSvYaQZuikyPQ1P3PqC2+mQ6/8lMME58ZINDtgMbo1ezlUKL1rWu4lCqUHtP9/s
Dj777Ob9pXT0pmDieEyygNH24IQyw3Oc3chgQooCq/+NF7gfyIPDOJ4g+DNS3VrRhmf9Q3M90KXs
5UOnujvVp9g2vpJwggK5vcF2/81Dfo9d4EV0ONc1dh67bMopn9YrbkPxZ3FGvJ6ZtEThwYcezK8v
XSIJZAN30OsgqKg5DWYycDhb16E8H1rPsLVNO79XdZrcJhrqTyrLxBUJbfX4Hr2rAp3/UJVN6Ly2
fz8/vy4wFSIqMzNGjgdD+PTQQUCt6g/yzZAm2XfWaV8hWwRIdXlTzefd93Lap+5HnVBwNvp9DtjD
DNUSOBSqv211RqZBP2dqpCJqPgOP2MC/JteOKYkHMMieZF5zr/2O3xTqCRdH92Wfwiv+hWx/4moc
26enCPW2MrcyNuWKJnY6704kIN1wajxo4uSa3U8GKA8dkQnirVWYse4EAYbk0LFeqdiw8L5LWmoB
hdCrJ45tPS4qVqUzJObA0D46+6S51wO37gKOcVHlfy399I/wkCxU5a7jXXl96BN/OwKF1tnOhavH
bB9C77RPKH3YWLnxqoaw6Dilcg5qMDFYAotUkeDRmywfs2mWwVhvET113Xto3QcnDk7a9bc/5R8G
4YR9Yq7qshn9btOsSzXiYQiDjcswpvd7vewmnAwNYTsRAR9GpBc39mGuApYPJo7Tp60Qt4Dc+CvV
/0H2CEJoQ1UwoAZ1j15R65y8ZS4RcIl5CzlHo2SgKG0EcQEQlQiBhCOjmcOAd200jU+lQ/EqVvnx
tJYzZocRILGNJn/dEgt23XXcdLRPT+O1b016Ho0+nO0UzjjpVte/7W+q0OIAmW32Em3PKFsgqOdY
gfJDalS24rg+2Rj6xM4WjVFofvsrYgbkacDxMxY+OTBi4cIa6Xhzy8qIllK5NMbJ9hLw6cs42y5T
cWI4jtJpj2SbJd8oTjK2IWmaixj5xZENdTeAw4H2Ou7XhY+ElvuX993PZFK38UlvpSgGBbXWqFRc
571ckZI3fzV0sddsoafLOd+M+duKSZkI0fgwnMxAZwE5EdeGO+bhnel+/VT9jexVBMQpqHG/54LA
q3mtthwU5/+e6XXyUOayT3J20bOZQgUSHnBLxoIp4PSvA/iqWyC1Nxxwp14o80mVte0aUIN9+0QS
RgeWxGWioXCF39Mq24Z/q7VC4bpMtLUxFom1rvQn2FEjIQdGlyBVBj7scwNjtC1YXfmN0fwZECpa
x1BSfhmRk7cNRxN8G5Mv+Abdd2yXLdv5zGaffgYM2Cfi2O4tWLD1DxVM+sRV0yOlzjBwPhlGMyN4
HFgR8v0lxkUVJPxYMTd61bwKwgQ2wKxsWU9HsmBniOotccEEtetmq9oCd3Rr4kLqPts3GrMvDR8f
J5GvqBvJrJlBp/b30s0Jh+Ureo8HDWL/sfA1aeRq/v66ZVGRJb5EkLp6HjxI5Jbfs/wB9CdG5QPu
wiTS5J9WgQDHfFKVvQPXm020mrMSYTHDzahI8yY/SpoqQIDTXWy3YzYWkvMu7NnksvmBqQbA2rXA
nL7irIdOcgMlnZXwtIL7m71o0076SZ6vJY6d4cnja7zAy+cGEcQiXpCaLxuAKn1zlTpUg2Auz3nQ
wJuhvpXFRjkqudGMMT+ihfEd8iy6vJk8ZV3eaXIDCPiwntttYc4bET0nMWhGgCjq8yodej1eWDUS
m/gp5Kxg0my1LAcXySpWfxy+5CaKNUqWNUvhilgz4JWrIZLrPkB6Fcqnu4Si3Huf7RPI0eVT3QZ5
dFzyCuRdkrCn9BnA3UyfawaUcJpBsgodABSFCMVrBk1ZfNpDZVg/tfyF1NXeqfK2HZPHKZrZxRXG
Xr/GTNWPXqLW9L4MiMNNKRW3uOSLRPoaOVEsf0bPYncZtfC0Pcwz5kC5KeBUKL5Pg0oFqnlnmoiM
SnpbrS/wIsL/Mdo/hYsTlujeVW/LetCsi8nhQgHOy4NlBLS9R+BSQ2Cx4uvwpoKFAvlonL9MLdIQ
8sWnJbGzJxpSgCkQesKLTVevj9PCuZ1B7v+YBOq8+0LEkMKxwrZ5FuXEee+mrZeujqYlvCuL7HRL
uLRTUF4gn7WWrVkyXEBtX0GmEPCTlHHipu/lL0FyKyyw5Gt10Dayt5N6hD1ix3ofi2GjfkUHNTaD
bnW85ZGD0JU6wM5490UGLTIfz+qo9r2sUUHjjSB3snJzbP6ERbojMxYKa6g7chMON5MoNqTcUo6O
RevVCKEyJw32rgSufjAMr0IDSst1E8eaHZOmBdZW9mbLbl6DQMXIWOOX41BF2h/Dunqphv5RVoi+
2YwUqo3GNrV9WIIoyX2wzhL/F6u7o5+nlsbENRTjJJciW0smnPT33yjOMn8osKD4fdV/Eto6aHbV
I2CBsQyZI/e0EyB2e3NYT9d7Dl2R5d6QI9CpofH/3d/Worfpam6rb57sxj24yZzDYTKaPM/vz7Hp
Wk3+djhKMHaY7Gmss/OAzoztKTXo0m53UnY+OPq3MSbGxr8spf0keVNugOfbqi2yrWGu2d9+7wv0
ryPPx8H0YoDUfPEJ0L7X7OcaLpfR3A7dXFOSVFx4gcnjMmOfwtEyK0LzeMROphcgYhOZaqWmYpuS
4MqxiBwuvKAzufW+ca7efOqr0kt3UKKA3Hctgk7EpjdAaOnwTz+AvUxkW9vn/9v5vZao1K9ec72N
Ab286i0y0tHnTAqtfDJ/WGmmar4ytg/ErVEI6mdVd+4VjMmMkYDL4T03WrFg4PHSM2x81tHwli1l
OGnV7m3a/aLqbEdVTTj8UtkWWpwGm2ua5HdFPIEiXmUyRt4oMaqoZ8VgnjV6vTILTWdJSreGDNJ9
yXs2zujgNd+NxqtXS9Zinwv8pLQoaftwhClJUM2hBG80Gxchg6KEoTJmzfd9xP+ttDEIG1kCtjBw
K0bKzA3uQ+CFyN55nL0bBkFhcVjaO1fYP29EJ9ymR3pxG8/r/ZW+Lso39PqKuphSZYqmzvCM+4qy
9M/rwApK3117YiFWOepdnRi2ELwSY0W6r6f7zISMM6D/6hfLglAePXkRIdE71WlrVrnnfqcJUWbB
MiW/WwD1a316eR3Oq8njVXBW5JApXWL2QUSyUTWXAruGPRH1CbSCCGzgfvLF9PP4Xg5vyyHBjtoC
4eNlfs/wAzycK7jjaBx2dfhW+zlyqgtpeevkrGpp6L9uEDJtvePnmztloo4qsz8S4OUKHLuR/LN4
2t2JoK1glpDw53YKfjcaROOw/ckGCzw75ttA7RNFZceGwNmro1ikvfO5ePYD5ZfB7OEHy8WIl4r0
t84krLDvHOVfzqXu2rVGBovtzHdDRZJVhYdDuD3MHCnkGIjDh3h8jG8PyJC9SYvU8wdINeGxYT7I
JyspkadSfQLlsUxNtNUOjjMxnXkiIDLCyUqRAR2+xqkfm4ibXlo/RC8z/kTvjO6GiByFwI+Srn3H
AbF77g3tqxPilQY7zkIl0rKx0LUbepYqdGhghP7WUSU3KBvk9vnCOJcoiOsvzxm/swX357QEkukq
K7v/ud5bWjlo/j61tSd5Zoi2fR14dn1mUeAgcXBm8sYkKiRojqnttvFkHKLMHkLuLI5c4zxcUj3i
kUhSHCWjTvfHtM/G2eJEJYyvvpVrzHEo7Aqkq0G+kB0BHeK16r3Y036UPu3vzWuWW+4gOZvO+em0
2/kPj5H16JMYN94QCUOBGm3RBboHqWWIx+WqJdz+hkpXtz+4T0AGUcwUh553pRjl09duNdo0eClz
5ZWCUO0YsbqKCeMZro0MV52/YxHO7rkdAbpdwunWuSpQmEGkvjOwtC8RO01vDKLvAYQPOXhIeMei
+QOZvKi21VhuWvY+qm08H4/QMCzGKbPgsPBo0Dg3NwvdTyjqLVA8RZ6GpVEGsrLG9Clrk+x+Zcx+
4jF2bpGqgewja0D9FWXurO5d3Qv1ABWMuV+hHvDeBmyRAiBWI1GTNsrtnGl71GvFNliUl23Y/wGc
xMcsnUILdNw172DS4XIlgSzB5A7PZmPOG9nd4iwGJ5J8L+2Y4iO/jUlQSzYiuOMhgPFsgUniIW/f
aWzxp7fR9NHQpg0o/qWfYlYQ4CA6xZguhJXJvWrz0YNLY8KqdUzTGEUaxp3WAhzCXEGqL3nvTVIM
sUXgxuNI88eq5wI4IoKTSIUcpRbi6wJ89zIe2N3mWQ4CZOGyi+IgfJr53ewmvMXsZSt/KpxnPCCO
gwZ2Absx2m5GyZ/7JuVOErK04KD+gWcMGQ4cSQ50gk93kKrex+MwxDaFhk0GvLrFa/L9ntZ9wZ5X
BMWoJrr2SXSRdMV2ZmfWZ7YQpLRfMuNvYXf2Sgcu5sndoNrORttA8JYw9Q2WJES1K7b6DV5WGj0O
isPfPsZ3lvkfWNeV+zsd091jcbgZWZs9GHH10KqtN2JIlGFWtRMsLyYNKZt2eZWf8pjX9PIF3aCm
Nk8+/LSqKBxQd94WHXJQej+6acMcztBADUQDNR7n71cip0ypvTu2Cifw0OPM7wLiYRnpVOkhKgPl
ktv2tAdl3V4ovZYXFUBz8cX74SaFbsptSBPC/1eqPRaO7Gt8mAEABVxkHPp1+B5bw6K8emGHPPlZ
S4S0NoAbaVyIGi5bo7I57FSA013eKxNJtZFmkyOpUYAGTXu6eJ++d0ieKwtv/iA3UgcDrJPEe4mA
v2weYOpfX0QiUTSYZebnqGIh2W9Sor6v+8A2+9y7tBHduPH/vjYdxHyyzx741w5tz6LUnKddu7+y
gDyg4LQKsOLFHqLmiTAHQG83js9MCXRuXQozPry96HXXjoaWqCD7FJNtHB7vMX6OxWoz9Om/Og0I
d+OmE1Gbk0s07jdO7osFyi4D0oimInXC9msbz0XGxTR2yPbucoQOcRihj0eiGhdHuvR+UR0mfeAY
urzWanbn4+fFIgzEv+GFW2/Zfx38eLnMyO01J6P72tHAq21XkUt/sXclnNeARzklwuHfO3oi0tsu
q9OY24LehNlQt70vN/D+dze7IJuikY4adGZvAONnuUWMU6PYObgLul+zkUi2+hT26V0hrv/i95rl
E7vIHySX1lZs9a/40//zw+4HTrpk0cgIRLpa6xX75udUWr8+WUYTkv3GNAWvLFrrLKbTM+l1OwmZ
AcRlXe6noB97W4oJYKxKFaJPLQVKkruVNu7Ee6DsFxvHvSfJZsCav+4RRF8U23l76HnpYZlPNg9p
X7XUUaZ/pEiB/OmQlSCuer6dXIaY9oxSS+L/AUQ7h+72DkHi4PsejhogShh9PrCkyGzkSrUWZprD
4Pv032l1QPJ6/V15t5wbgJy+LIVHUD+Q3RxalBL4FDy2QLOA119e+T47NSWukQe72RdWVgsnOy1X
HNdNm0lnuDnNL015uc47XEkrF+65XMjgVAdaiDFd0Axp2p5K2c1HpuL7L5ECwaMlcqDZ6l9/8A3R
eNZuAUBpNcBc2OJJnXucmGPM92TU6YDrJ4aIL7Luh0+gHIilRO4CQtux5faPxzh8AmROqgiEACw6
BaAyEXOAr8LFDhHYCXNAihRgDU8iBat0Btj3ZQvCq+cZZK4qri0Y6FI4pebJWYnmqefa/b4M+8pa
6OcvWy3lk+UnNOkNnI70PXDl0ELatBhPA2ADeIQGHogkE7NZkgT3pGLW1IAieu3fNWdHvg+rcXLj
jTd68NWqVKTwOegaGAZjXJsolz3rF26GMqKC5T16uf72BjEobi3z5lG4XvIqe6B88gELxKeK7QVT
BaRAsfQrzw3BnHBk21A2dLTs1gdl/Xls4Mc2ig4Xqq/6IDmbXSKiR4BRA3d/yLSs95yKW8dujZ7k
zUi/p2nF+AEP1nKlREZXl7st2dmhz3Ubxefspdb8UzXuHPNradAJMXvw65Y9KR64rxiYuXpOEoWf
S1+wJcOS5CKPsG9hctIgHvNS2t44YwK9YeC3hXx98DGHHNUm267FoCMwuA2VIWYx1TfFPYGsMbWY
pLzzvkgSI211ZVobH4A5E9/G9M3cQqZg7aqcco/f/x0glxIz2gp5clr2jZIBc53julwa5tO9No5V
3lhbzACYJtLIDNJElSi3CGNzInLSMN+teg1bvn8j5ep0V05JHLBq1v63KyN+7sArzfa54sfLjhnb
aM9KsuqqsZjb6Sx5LkE6k5AYr/oV2IzW4pZrHNohaBVRKbewHtPWH5h6WvMi7G4BIqSbtIjlckr4
6HLAg6m+058Qsrk60oiLuFvARLetY3OZZ/+jNkwojCyrnDJApdrADdNuHRqSQ0vXB6F4fMlfLZ43
2gDEtelbbY7Gh1DVK+syUP+WmnE4ow33ATTeTXPCzLoW53nfN+x9vanQMJGGqlo8tmqLojWi4VJK
mOn1caZ/s9rUoa0QuKsYrA9jPYAcQ60u+XGYftBUEM5F/5BL1z+Z+XSFmXUMH2u4qSdAFo4WHQeI
8k7qXcOO2jpSFhZpUB2tmMldM4df6NwSYOgvXubOBMqVya/lYhAxtvVuohsMXkLFeIbmupAwmw1o
XY0vWNhzOJzTAh88WlBtOKsH47GoIOw92DeIrWpNlj25GICxHLIPisLo+5FEePaUK/jU+8F2GD76
RLgl4b7r0PCbAX3OxXjoX2r7SuvZjYcicsAMXpGfgc3h+cD1MvezgFrCQPjN5HiD6CUNRSGK39dr
RFmhJHUIpHUjQh107SBD2Fv1U5NnC73PHIjjSFbmpP4/LiInd1ZtuT8x42cOsT4RNWFl/Ln1TEix
4et/AapLgEGk7M4zLKWYD7bVVpzqf+tR/PKLH7NWcn49NiiZ2hRHMQmTPHgWiY4xioQZsRPqYmPy
Cc6z34d9lqL5ED9a6baY+yuQgoh0MzsxnrEPvOufKnGirsJu4Lww0L8dAiTlbEtRLVYQRGogz35V
3g8hGECT8+Z/bB5xBzqLWZhYlvmiwT1G0hg3szVitC3YWyL97VvU4xO5gNbKb+6KcBtxOU2IybRp
qA7vgh5Jg6TFMnOcXJeHyLtYylCRROjvHSGH4PgqUAeCfEAPHBtu4F4LXuLXXKwPybma2sEVaril
jo8DVx3r1sXqGfK3/iMipeTwrBkNRIqqq86AMqY6v+uyjVfkrCqlMKZePlcwsfSVuulvFJpSfd5+
fmowrlacWN8cjrdmdVy7CNbDTxyCZ+XivxMz/ONAneVfFyZqqwGcf5Bq1DR6B44bMFr+LBaK3Zpu
xHYnu1jN0ogl8rfZoaq8rxqD/CZBFb0cYVk4quCr6oVMJ5TXCrV2eP/A+IJkmQEF9Qtv8fbO+hve
oKoEjTNmh04unZhPkkkOlTY6z7E69RTKAXvVOdgm6ge66QVjMJVS+RQzBbak0UOTXJi/2FGDg+Qo
O5gLHm/Ums+CVJEvcvOVOuWb+cpyhfTy6jJEgmn8yZxCO3MIPp/QqIQALuJTgCwtwuClRz0itUyd
3x6Y9X6EbhQKYIpcHfr98U8eFim4NDsAJe1XdlwKJSJ5t66CUEGWraYLoCx/2eN5x6Mr0SU8Our3
+TqAObE80JnhGQiyR59XPHYliPDgDe25dMgLNxiy5w9ONL2QNa8tqiQRjYtLTQdPEZVrWVV1oWHE
/ySdrJFKL6d4BckJEvY85c1toZ6lFbrBO5oQeiVsQ8+PmABYwNRJmLyDBtuDw23/+HPKb4Brarzl
K36oMocbDg50Ydg8pMOkf/CmIDmup5Nd+hym3nmKWCtazyfG6RcjdfE7baideseOAADGGPThsWPU
EUMS9jb/wYIDsEwOUWQxeERfUl9hv4MSxJ2c4ZjyHkb6ewwZKFYNTk/FlEiS/+W6KHoYJSJKm9Ys
jtbZFkiswREeWYiqrODqyyVk8y9Yp0uUpo/RKJn0LY/a+RMbbuFfjF7kQ7sDaoOb/Z7dsZj3234p
z4IOK16Dd+OESbs/WB5AnZtHwgZ5pJ4dysiRBtQaqFIhPYO+VmqfCBYeDLkF2N2tqKnAHM6+8FXP
wkWUypHwbAAZpMqHcV3MyoKpG00VvNA9HBTf7JmMXAJkV0Cz7983D2130vNkS/p4eU14aaQ6bulU
Bpb8w2RHidny2c8JBzM4IB1DiN7yfGkXzSQ2zOiNHte3UYKwWCCr9cuE/42sSNgVACJoNvxqp6W5
z27CRTSFGrhE1B5BFIKKZK0Z0PXGHAAPOmPz6hsaTxOikUZp4ZGBDWA73Vjeu9t+ebvY0E2UtGn0
OVj9E6k2FJSzP5PgcpGd0zQ/xX8+3AUNL2H09o7uORpip6mK7WE/ZpO4DLxbWXjc6WIucTNNijrg
SkYakvkGhn6auERoQhw6VI4lCZRyiLCCDD1H2mWevRUZ6WxKmBeRLRAyXDmGEgHLvoiFk5wSvklY
uBM1DFPuM0tqIhqsSmK9mQs0E6W2vUWZPvOVy41dJdqJ2Cm3d1Ifpqj7anPM5/2byAKGLQD7pTwk
IhYadPDgRy0IywJ1R+YvhpCDOmyJr+bBNw8VEhQlR8RtOPoeEnd4XM3lhCrotbIh1n7q8Xqqa8f9
hlYlOCVy0JDIDNphdtiUmz2s71VY43PVva7lEsKfN5j5A2h5sbKby3KT5Z37Ze7s+Riou3bIZ20j
7jlTh9zbacEeNbz2ZhghDr0wAZoDuqqWeo4hHbimfHV/J9ZZabthB5yeOm+liSOW8UcqvHkRZCeW
uexza+Cm7yrzqlYdQ6Z8IOPVxogzcwDp14V2KJWdmFRpMTbJa2wd5tTXPeXzAfwv3QIujJnookFG
nQm0pl5ptLMv1mImN9+bLGTrYuQ3RLS9E4LmUG23n0b1gTH0C6O0293EYDFIipjcXPzKnd6IaBju
RwgZyjbd/bie9dlA4y2IZJFAFToTclyng+Bvnnp/Sqs+lYCiYFs069UkRG2E1lix82jfCZg7R8hp
u/hLKsCqU17cXuk56cCiXjedVvVWADHRWXskp0QViUpl4OToxsanJpt5VPPj/FHzM5hyS/fGwGNt
juOfIfD9ybLp78kwA3KgwxEKYTqRW/qLSTGYyhhv8TJqEi4Kq8U+Vc3n4mH8YrtItAUROzGq6Bwl
/ryqqghZnLyu433o9m8W9XsjVygysBEEEPOirsayNIMl38rnZf4t9HpDZrf/m4oJKoXIWj0+Ya4k
iah/zJybqboDXqHZ02PzABo1Nuj4l9CBLWgeWYbJxilkumGvHOalJ4MXGqM1O+mJwTy3VSbQTxet
Zb+jjkm3/5qvvm3mkgczcT37QQSKjBGYMGwaWFbqrzPcNftIlqKBh344QlCx2/EtIP3koa772SAq
Ssx66ZgAmHHxWZWM8PkDwLxLYhx1pKHhwNegOPZrlZbG+rBGBtRKPI90K8vpMRGxaheSM9wayt9d
M9wyb2JIpUWTnBNpml5Y7ubf+wb1lhI8R5EVHemnxjLYkoZXyfdk4v+Ohum5hsUYY+E+/fiBX5XG
Sfgdexpokn9s2lR8owBg4CdER0DI2NbZ/2b2nNu9cONrzVE/iSur3TXHcpfj6oKax/MSHqjf3I5+
gjlV/Bn1p363+5D/SnZ0JBnLT2ynYGky79gz5TWvyU60ohqzaA/rTdVN7cgFPxqEsKjYq/xHfIXu
z9UVvJiacz6n7xAWEg20ImXCOlYRPbuS1+V6vcHyNPSN+UxONT+2FDGreMaIL0JCeJLF/S5QU+xm
Ing2K7DRlvasCw8Fm7yxk3vlqBkyLn4eBxfQUmI2xamVTxSKusZeGA0TA7VAOIq/2ATPAzwKDSuQ
9ChrJfx/UB+KrV+HvPrBaDit8PH5y9+hSimZdCv9SP7kSObC+2HPgXBN+dmaL6o1afAxuJgMqZ4J
CZYFUOTK8zDmVow9AOgBswUczDtBDV89rO2ReB9mgmHgXi3ikQiX7uIT1LFuKsnvNF5fl8IJQHxf
mnO2nDa5cq3AggVkzUb/4ealVZD3w9WZARncAVFwE7cGXpztWbcUTm1XDf9jKRy4dML5p2yMPmVT
NBKO1+d/2o/6IDeMdeD8nUzdgb/wItQMFIBCxahVw05D0tmSst8dOocJCdvJdkNVFyuR10k8O8AE
dKE1nJLaQK5+4wGeTZ5G9sIK9H7hb0+hhZJCkDsyKzgXbryhAVAnPFY8P3LJw+4saBmvqqq2ZhBs
ns84N9G68s9CPjmvbjyPHsXVhfLvsmhQ9Li1srdCwvNGACqDRXuwTaimctPv45uEMOYiQx5p4xy6
M8Dt88r6//YCe8GTpKXt5NURV+upcSZDzPe7h/645VR9x162gg7AZ/YLi3YWafgkFaKOseSD7pEp
kg7izez+NbWdW/HqcKVNXsEWEIKe1UPbaU6mX/S/yDsMLNFIpM+Kj2OjkV8G7vbl5FoI6cosRDrR
+qM55EC7lkNi3anUAioCLE1LwWLooeqkhGLoVMMe4hNYDNTPzeakc+TwP1brptnfOfHRTR1m4SOQ
4gT3bhijAKKGk3M5p/OxQ9l4rcSWvFkNPU8Fb6ERInyzbY4Z+mWUjlKP8mMUCtLJqy2CJY4p3j6i
AACb2Cimv7d6hy1eLOW0LNR+G00BkVLSpPAnn1Wpy1ikc915BjeypZO5Szss8j5IZ3o6YtCcAfkm
bJs1UWE6SwbufQNRE/CorKs2XxtQQCHDG9lRbW4/qEcqovcNlqq3bW27xPfmGprwcQiQTM4y7Gvw
O11ZXprDvarZRa7ZvFg7GHAa9jXJPbSd95wOz2Z/FaTDVrLP3JGBOlbmocCIkcruteSi7/MTsuRv
DKigK2xbZ6/I7gni4OY7ITxDQ7r0YTE3pw+ju3N+5AL1Jd++aHg6z82Od3yNwuDhUupHKvfcnoEn
bIGX+Lp9ieKOCAd5WkPlYS7d+pI8XS+lxvW8RE2SPKkDC5pInukWeSke7K+1RHp048PoVNHzBVbj
rYqLwgYCHTeQlGI2ENVzF1IOAC3ZdIqvJ5h7pmFZmrgMQohal0SugZ42lSeuTlCOR6Nj+InsCKzE
hip78HopLn5t9Q4lkIOxs6ju8V9fgm8o1N4QddQAaM9/t4IBvgOsjBEKkVUaWCPzGjvwzVsr7qPf
WpxJV/33yYZpIK1Eo6L7hb1S4BTCs0mdKmEzCPF0XgLPEO5H24SLNyAhFTsUIyGwBEBY63R30txj
d8QfrqtvFN4uXW22Js+e5BoOwT0EbHz9B0zqUmUH1UAEgZ6CaauKwaXSS361Fc51nty35PLK+W5J
198aNuUAxhfOjWOgCX0Y1KKgmHscU0yg3XZeOFsEawudhUn3YIovWGhoRsdVU0X4fqSyOFChL7+2
F8lMbjC5qVmAcNmcGIZAPkrDyJF69LdmqQeIIs1MoTQTh85tq7OL5+rT8x7ZliJt8ywJXaRLq/Cu
x57kiwBQUZ3i+4daBUkIna5u2GfSb4qdrjXALruaWNCBWxj1hafB7DqbYyDqH0NVUk2dYfXtmuug
i53qSYJU1pQvo+M0qqrwiP/Rlk+eS6R37LePtEXl0NGEvt/O7ZAFnKnVR7m1W5WWQISZLBYK9ZxG
5g7OqxGQoxPTsMcheny/KSt3ulEM2nHVEcRaMMq1tYBMmFjW8vSit5iKTKpVdE3fV//tts2CJGCP
Ql+apWQGDiCR9RlgW0Drbr9Egxi3zQH1SEcf8rEDCl3bAec1Zs0YRjuHjMuyFd37FCDVz4HHB5jJ
4sM36wWkeUN5d2nsC+Ffca+8wbk4zDPX23k8Lykp0owizCoDd68NxKoB0clCxRVjxBC6sf8SOwsa
wjNQb7+vKb/lkaFod+aEFRc9v3OkFPwAC52EQBx2DQ9WkypI3CJ6sRNTXTDUw931YkA9O7+PgFT1
4+iPoYNbeWCpVrYmaOMVtQTLp2Y5u+QZmOpLkBRtENmEkbt5JzFx5hCNkNwHgwVgzfqyKazxi3Uc
0hmjkkwgwUB2f7SSpEDfcRGvxF/2MZLFgHQhaPZpHOqq3FISkhC4GU8oWBXTAnW8tTK9zEOdnlz4
WtTJvafFV6IBxWOZMp9BtJtXO5k+ooueCfpUQxqFn6tZ4Vpr4GDXBClCxrgtYOmJ/wqIZg74rKrg
1tSZQsiwykAqYQvaGJmSdgsjELcI7iko/Ycn8wSPVMsHfMrQvjaVpW+EWV0jjV1pTmNuXNnyYuId
LakcVg0fLEqiR86fgwPvpO/ld2Z4+N7S0Lj8uGu62vCkfF267Ixu4HzFfs1MsIzyXMfO9CUekT9o
8c6vnG0YAbAV4A7pGSzadW127Eg1eEKIz83pPSFrgS9IeQgYUGuuIhB8a6bJ+vsgE7KxiGZGfo2h
DlaFcqy88i7LyLLvLZzOybfXlrIGZFe3lJf9QGhFnbIw/XwpwvG7+TMhiqyYTSgeFXsOUFu7zUZa
9mtjszpQoWasVQFCUf7N/TNQugUJm/uGKDFO+ncEUAVWtrDBF8naZFIwWNOkAPXUsbyQ6GnrYIIw
KToF2aN/SRK5T62zkKnl5c1EwuBwchA17fpLyxX87zWEyb9y0E5Q4t5BqeHZ9MTNibWR2X6AUZu4
30zHRCxaEESfHrbkbzXB8nfTgYDg5fah29/ISngkbFexf5YUjmyggsig/Zn9ozqjIwmIe7GHrCH6
lgyzNfLnGodXPY6IHqCWBl40zTxZfuFV+GZT6GLLb5QeQ1bRpvZ9cRZIcngj6XGF57h6Dilt/9om
POgxd0cWsjxsdFp4MEQwp5Lt6ubBU3FB8TR7MjL9DR9XWfaeDXA8Qgcg0YgAXK34n9FdpdFc4OYM
QQksx6qp+RX2Lzj0rDP7ypOC6NWeKiWsl+ac4ZQHz3M1QfMlYTV8z0/eqgk0eIQcOK14t1hKy+K3
jIx/NrLke8YKohW87BU4TV64qjsQ+6EZBmoiacb5FKQ09xZw5y+4pl9iqz1gUZzZfKAGT6cjQ/w6
mO9+VRIEK8olV3mMGOTiLWldF4yjZilgURgxhpirriLyDexnJQrPsYUrvSQTiQXKYVRinQqnJNp+
ORtLIv4uQvb6uDFuF258prleoSeyTeyGlMmJDMyWxP1BCdN85fA9Hsmgh/9/mlo2oLkxQHxw6DKp
2iMm9kOhqCUXIrjyzAfYQNT5+EFg9goD6UCrCF+amAOq5dbh/On+HN0wlKCUDRf2qwRTbVPO83Zr
3Y/iWlsD+LNDqczX2UFDzd8JTGBSUk0xzceKH3fQo78pu+HWSVl0yAktIc0rPGQ6wLk24WX017Kq
+tFzl0Js3J96OmOwyD9VSD/a1XldPAJXPzI2CFxJZRGG45HtHK6rkea8DuECix0WHzky1pXmDTOe
J0zwxhbXuMkY7yREwm0+jw89g9v0T7lFJ61KNy/Z6llHB1/iEKik531xA17+pCm+n59bkwV8Wfq1
INrk5sdTks1UlDhfpT77MhGexOl8DenPl2sZgRWWoftvUXbvI/jqFozhz0Gc9MJhsknk4B3ZzAtK
0QXvGhkPeLJhmB1sZjw+chUaMc1+2QaFx8eBRkvHx2Hhb6SOvL/qsykPmI9UTIQnNL8yctwiZNBg
HKnxrhVDdRR0vI78cUk97HFuuLj7fcVBdN1tC+8r7k79lwGbjkVjAC9+2E/CpIIlSGOFaovVdag/
/na4pZ3R34e96pcnPeXah66adWiGpxqQ8gU0DOezEDlIc5jwHm5z7xJZhTpLWk1WOeBNN7LUPSkX
NoZEC4EmGcQjf5ouq9Z8mXvqlfLJgfPLEnc7tf16P6M9ixwB3I83jvMBFe9aLHyEmnAfj/iLEoyg
+YLwSXmSSuaRhxMt299arbYSaGDGuw7CRtoPIOJA1UW8/cWt+WComZZfHVuZLsxtRcA/1+BzGLmd
Q5kiWuK4gzUd3HhKZsRow6t3ew4VHuhmdjvS7BQJtU03gyQNi64d7tWk5aYyUEtsykhqxRu6wgHl
OSQkMTve1SCiVvSTUFr3KJCgUanuOl6rSr7lYXfX7Ltv0Nvj99aDGCGNnA7f9lcgnW+/XKh+NqmX
m4q+6wTK3/NSukBUy70mt5AxQ8L3PxRy0LiAyUcFA0ifBcRZf3DbTYVHOsFvLpWx1GUlwMu7HvVq
sIWVyzBlKQdxK1rXEry2Eiqz8+zr3sd5HetFaKbEuR4KICQ36K5CIjQcZt+JthUN2Wp2sCU1/iOg
gl+2OxWVJ+cadIl/b021XmicwE+wDcYkbcmSCo0uvHCWob1on4nYZZ+rdkLgMac3guK7YZQbdpdm
uIF1/J9g632Z4u73qI9JBJjuLXBtY3zha082onCNGPxQXDwbqxG70pQW3vQuY87oKPIRqvYVoYNE
fuX0vokGqhAA7+cI+nfC3IXtp2Ecl7truyzj7ADTJ23pAtSfXZ0MlvN1iWArlzbFRfp1KEpUt9Ml
OsGao/ARyHnOi74KF8B6rl/sKwtEtoFKvZPifDXtB0T2etQjDIBikpuxMjlcyc8qMB7XxTCByfnm
H1+1Flc3apx/B2Dh5vc+S2pPT7rV87c8X4ND71DzyesNGEvJFycXELwQfBFZgm4MUwpYEiQm3OyG
01Reu6623O69UwNs0PHK8e2mRRZi8uEaJkIR0LbC54uleNu2UFWie44iyJYE8x5P1Gpnzrs0n1vo
Zs+WK1FuktRmdYPtovOAe+jtzTwqptilos0Y1lbSimyQPW2o5VeAQSqvL6MkdcxXquOGtGHGyh65
TNiPNXQyEaUCmcSsVCsuA+zlTz3oYkUfADY4VU3IT76g2TOLQbjAzazli/cIqQCrsf05T8udLGpO
JsMLxOYZcZpEoHXkWm2AC4BB5f/XUU4VwcsCdTCZpOrnrJtgx3Tcf/+Y86zCwXFzncgV1Ob55iGv
mBRow2ADt/c7EjoKlhqjCtrUpRSUTAu/VV4sIE4RbEI/RKEqkMYKUgA2JhLkCUiHxAAFtsIUAZzz
YIVt0l3mNurFYuqPd6iGOaNIKAlTk4BcsJelPm1JYJZX0RAsgmoM+2KaNlNVi6OPtMeHJ511dIsZ
3hq/QtPmCCGjOWkWFKTDqyjPtYZ2+RpAnTimzhIh2AWrqMQnf83diUBce/nyBh8cECpF0fSghLwV
42aL8ewCZZslrj6Ee/1F4oE67jqhp4EwoUSV3jaezrvd4SWZAWPaP15QXgXuES1OowZIPGhOq+3S
u2G0t0YVy/JxKrVfXOS3X5P5N7vvcKNOrtNd2c4cKmjXxX2goSoMRczWpSqvRF1heOKS4ucU/s12
080JB1jSK1oXjT/vNoj1qzPRpJ9itGDQkrIYLSPnxRq19Hr7eQg2iwqjC7EAyjYNPcWp8LAaOGJi
/OPZUB1K9p3X0WHkpSgGtRve9grZH+Di+KMmpBHywIpyE9HeczByRGHFTKIm5fMdsoNKL2HTub4V
tvQowWRQ9lWNUm7BC02atfcIb5/NkucCZ8cT+HI4YiwcgSkZ7xLcf3IjHA704rFnO/1N2aIpBq+o
Ano7eQzaGNf3tTRgUrf+HM6h+0ZRKkPrc5W16rfG1Dioz6Ll0kmELEi+ksaHnv2J97gvJVmv9kUR
ZxgLKm1ZJ+0A2RDEWKrRD479aF3GwCxb5wR6f3uuR05Dy4Eo9NUAisqzfZ93NMyinHaRdOFv91iE
Nxfcy109d/5ByHjLHlcZJkQCJfKW0sOjYjOZLFDfFVpExw/ml4xf7E8uFl1QupzvRvMLjYrUUrU4
biNxvTCffcqgYxmJ02zA54OXxudAQl/HFV39YArXyu+8J14H2iLwskn3SKVVXB3XoBRvYdaEFAxT
RYw0UCbsajpx1usxyQA8A6T7doVbI3Z2zlt2ex0fAK5N1pNbsxxYVQF1+2EoViNrczupv51115gq
MZfflT16vspXF+NiWLjTrbak6nzZLyR/zrgtMI9/h7u6MvrNjUpnwscjnzmOfViDaQbunThRSh5R
R8oD4gAK+IudXtz6AVCs5kSM9TUbXsqd2eeXsat5hCNP/eXpzf5mkeTtunID8s51YvQ1T3AtDMGV
FKR6B2RSnpx70/qH8SIj8CCNTkXLfbaL2crLw6Ee67Z8+q9XjhnLoz3tYslS4Hr/HShe/hFD4Zz4
gZ6ah7oTuuR7UHONy+eNSUQbwJg0r/ftlzPiPBfxK17iupKnwFQZO7rGbnnT7wEV1NRHUlKgVdub
E9NhVjEzy/pDP9chFX4S4pHO46NTZEaFP1LJ9xlqD0Bm4nkleVc/BH13FA1PVQdqvaFVtf1kY2bt
yz0GJRykqKBrZmjkFUVBI+b+qt129xO1OtygKoiawxynxvFbgqxXpc1SVQo5a1XdYh3ILV4ePS3Z
uV1enquiHadHj1xO5Mf9LR49H6gHIFYwk2j0oWU10dFuY7OJY0XVqLcGCID4owfzIraCnm9NSs08
1nCAVEbVQK7HEW2as8nxevPHRYJhpbc6NvA6mqGgoquw0hhE3CQD5RVuI0yWq5izNYkc403klQje
ejVhwTY6NTb0CH/FEGyyteKyDKoVvTHzWacccxddmM2q+0CoqxhqUF+kzpvY50opjvSx3FUvDWTl
Sf04+BUPR2i7o2PMZsT0on5oQIiCyyBU0ZqMtlA9WD3JYayC71ukZh4pk8FAf1GU62ej/URN1+ci
qC0odztjfbZ+zXhKTsAWk+LhnpRiNa6xSUq5l7ql4nUztAUkdhzAd/3hpR+x2x9YfPrid1+diP0q
F6d1WV9dLWPJFyxcCC3K4TX6Iy+9fUlU4YYYqRcNoC6HWFf7pVck11JF41KVB+HDAHGTbNpng9NH
pawdZULVvDnlbs0efWHuQ8drTAjez0fLpGKsECdWnTHYMSOmRuSqRYfwoDfU/4oA2TjdfkB4M9Mn
THJb27wPv3sxFMj3UfCWoBmyqo1vz3ySqlKanNZjhcD9h/OtXb/xm1bk/pJsA65NA7VYVQfpmKSj
JnG0mg4G80Rn9Le3ZZ2ZthuxeBGqqesuLfOq9+ZJmYFJ+4MTNH5bgitzchkiEm32UyiUY6hE/saq
/R8qxjHL4oOOF9xh1nlsv6KW+bpMld+djqHYfAosTYd6t/NfAZMY+Qx+fFH3F1DUXLNl0SY9yTcB
k58bLlc2EWAd25P3HyaytTsCW9Ipze0xYLDtyb5l4TnuHke5YQswrSfczuTQPjE1t8NUPhoQjH3o
j0dgcwItILUo5il5sWRiC5Exq2k1/JdFPelR4zfVm93abmYQHI2tzmsz+0grcxbkfi2X3gQyqhlj
Jv0wb7nvp6ochAwbV/jzsi79ew6lrItIOVA2PnLJHlQOJolleSgXjGSskz3wEbIWd8qpdjEsSC2o
0lSjuE75TNz2rtwnOSGrcMJYN6oPEQY5mvlyVDqyQCpUpxRgiqJO3w25zcvABZwtKB56KccwqKuW
7Ci8PzjDwvWwEZqtftBQbPBk6S/KoJ/UTKYyv3/x1mdJsCbuhMiVbip+nn2zuqQIXyKOoph0vd8a
y3Tp9BBiduqb1BvsDmg3H4TRbFimO13K25oy8m3cSkkVgzbo3L9wU97tORbc2hOBKYrB3yV0uMDm
bOnTTGzsX+lICYZE53oL0YJW3jzpuUYDR+iG0BIJlhnGDTQNIVxCz/MHNhEJL5Y5R6I46AEOlbly
y2EydRy65GRMSZ+FwNKE7rrPaqRvM0jdev1kjFYRWF2hWni4qX0tAGe1PkEyKkgbcxbYFMhm16r0
IEHwVp+wTJNUPUvTT6FL2inCcmnijjzhDhY+9GC6HWGmvX/xNnugHfW5BHZpgXa7awb/mvGi2NSa
buKIJ/0CEEWW8D3z4HV5WSyY0rxnj0rVdvZ1kOquSR7NIrshUdIESdQEh7Rskc5+5/e2MOgSw4Ym
MGdhVvSnadHDJAFwKMsUawm09F6DA18Hd/5nuxXMwndo+f2Tom1xJN3tAoL0Ln+v9q45NCgSJtfO
Jr6px2V2rNgHiI2QZN34OLCnYb7Ja/SKUEQrFBFkaOjgPrFGnBs3VKQ0JwsZDe9WgOBNQlpEkiAy
pLG/yI+UFiUr7FXnvSPTCCZkpq5Q4D5oF/UxKgn+HO9p+cxipCZEDX7ZFEr14FzHyvNvj0i+//P3
LYrXukiNWFW3TPnQAlhgCDf2RansAtCkxM6VTWJ4YNQUKvjaCowL6DRmqcjALsbV1imeAfUX8oZA
VN3+oEmPIOc/BfqnwF4h1VspxkqSG7s7oooj4gYgjQY3co8S9MtrbZSlOK7gk0H6tEmZMtrKAHps
tWqTZOrBKPgwO3eDuFBTlFtr5p6rtpklmuXFXK/gbHe2xWaiPsEJRJ6yW6nDwZUAqS0648umemp+
01Id6MCKEhex+wkBAHzEt4Ee9Y9uGLFymZF6dLtylhpaNjZXrxUKxgpiwcT2nncOYHVDAjJFc2+v
JB8EdSLozfl/uTJxw3+WIqXFqWrfn4NAMqFhqByfXKXYUAyE8xEFPy+WefUGSZD/vBAXC2t8Hman
YfCtpvjGCsKJZm3X8B2e8svaeEf6Y9S5W1prP8CgwCIQKmtBmy5LUtqOXNxec4zg7QOt8h0J37SQ
7wtY+nM6WpsqO7ebN6cP6TvqurukvcyyUKIyWdiDBW5bgjqYqm8quw/msS71EJyTJvvHwivkWck/
mbKYRKtl4AzdAbQuubjpGliQ66qiVH6nC9pQmUMamsvopMekRfg7zD5+tC23oAXe1yn2m27HM9ca
n0Yy58s+6IPt9/wAVm2qzlSC4qxTK4DfC7+2kgaeul7fH1dSv2yWwJM0T+0M46Vip7YXIzWJbuN0
3+bEISXTo+l/ByyKo5XnvZZwTyduSalKJGQC0QO5/F0/kaIyTS66lTPa99hElWCeboyMuV41XNCD
1oLm6MMol2hkPgZN5GwyGZ6IFQQlgpgUSIigQWFGraNqGv+ZLgqjuW24oDrqz1FcogIvB6q8sk2p
Rf8/HgBcm+zS3mBnm9tsZcEBRV2Mjdx6QyFsPSm/FVVYit+Yr5XfmUoFJ6ZE4rEB3dhBwM0ned3O
XcyXSbxSbVB/wnCA8xjPB+RuKji8eqs0lz0Cw/aj7H8eoJJ02Shn83LS6gZxZ72E03hX/xJU8eIM
Axb38kJP1kZrMzjga8FmeryXUUyc889QgrmoS6KBsiRBbulQO0k9FCqLY9btEkzWVBvxxY5Ov2ZJ
Wa4JK36ef4Ah03lzYV531+PdevE1OnzLgob93ty/MAnBhy+9kiHirSUeDH+G9MKFV41A8kPFpV9w
NOurjvaAsqhv3YOlqE6WSkCpEHnIYeL8YAqzhSuE80pe58mWL0IwdySepe7y7Nm9VyuxAoUM9570
IUZ4zXDz78m9bMBrYeamelYanNJKtpzC5LLiWMXfGz96Ao6VSnxXrehQxyfZhBkMW/j3UHqWjBmm
cFCgQpfhjYepSoxtjS+0oaLiTRC0bWje2H48AKnPtY/URBBz6WtDzoxITIqEKajRpVKElmdWgC+y
GHCvH0zvkpOw+r651JtjiadDiz65Osgv8FIeBfU0HNv83w/q5khR95oxq+EMM6T2VdHyzD35jODL
3vnRs9u2QqChLO19CafDhVnoNOai/XjZJ5WP/vsjTiuOK3YZJ8jcZOZXREZonEhXUddyiR/l16SZ
9DZztjLOGHY3p2kZfvmmAK9vusae3j7O5RttFhlvYGOLCXQ1ZrJb/TwEZFbCnZCQkr8fOq04xHzG
ZfjvDp59T9jT7OvmlAAFohJuiWQ71HQPg6z5LWGYRa5SK3+/3kxVZuRZR8vUSu04wFVhSytcv2jG
/XmedGBDfO1u3daBPJnY6wxRky411RWKjMhxaGn1R11rxA4Cog6W8atIaKyzr1XDa0LvYrDm/1aT
XZhOPMnOImlsLI1iCOMsNE6ABsoTRE7BoiiG+kvWXQvdatRHRvrq6rvv7Rq7N3Mx3uJkkDduJnwO
xlwToCALw0FnVRQb8N6voPTNpR0EVQwazdoW/vBtCDWk8VX/3oCE9GzFetZG4A0hQLFw1zIbW1Wk
foatvpv6swBfTliYL9oaoQCXLFV6n5k8y1ojbkc/cvCA27EOWcFg8pxUnjkb22Uf3dzyMNBji76z
T4gK8wzHQiqZhNTtdKpObngREhDVIVT4ExnVe76WfpzhZNPvoJNxdql16I0dlU0RvMfzCWpRCcrp
CY/Ua7ehwOnD+9PhGc54m7Vwo9Nf5Ky98I/5AS6EWpSDI6D4kHtfPZxhBqtQ3JtjmmuHraNsO0Nn
zXNkho11gLhrE5bqZSOTeqjimBvesz19Pcse+qnzrrQHSfmW4MRd62sXT1eDqeG+CaygJomN9Npk
PHkbeJUUR7xteEyal+YVReshC8nJ17yA3+ikR1WmbZ2ktFZ/XaPRhaNnvIvYAnTJTyifVudZWzgN
96Obaos4pcpIJfvg5S7lsp+GHdTkNFBjYQ6vvNdlhvqphKbQ0hCm9WPFA32ClQms9bty5tziW8kx
1J85pM30QzWIpKxfo36vSDpQzmaw+wE9SZzsqYgkSO8bw4JRZG4PCztc4EG8VLeL+HY3ESLF1jeC
ly1bWum9uY129YOTsT/P2X66CGxfrmQjuRgF2739Mh8lRCK/mfCcPmnreLH9mm+LcDs2S8qXjrso
g3fpyoKvi8chmRaWcagF3SK3QFIgoGwhxtoqc0p4TXNuw4xNcuKJi2DNn/KDptLGsAHPlt07bJqS
VlnSUWahNyNPCPUlV38uOZLGH7PG7WfGLqkL5kgSD/I4eBVntd3nQb+i8FbnJKMAe14p8PlFsZvF
r/pcFdh97ToYmu1iI8rSMw2uxZfT0HQPbYHWO48K7GSuiY+LJe4xOB5SHhcadHI1jE+TRxMpmZGa
988NfFigsWdST5HAdc71tE9TUyTjEjmB2fakTiDd0GGAmcIGBoDYXYBoWgFdP8MZLvLCEz1rBZHw
cROiMihZnOD7jwjFZ6XQE8iDfQQW5V4Ab3tW2l/NuJy9rSOld/Ki7m/yQ4J2uEaPcNxz2hudmM0o
v91iC5IxMNfkeCKQSW/A915UJNmxuSVy4GitKdOvInT3EWZAzM1UEQoZBJqNUBFAFZMiX5/bTI28
nLZDAxi6xJiIBTz7CQwhoxjyCno06FVKgtOTE/Wu0Dk9Yg0Lps6kwikRR+KEUKaABuvlrHi/l/9/
F1NdgHJqiOG6KC2wbfpcXzCk34S7p8itpFrGngff0YQvruGKO41aSyXxi9z9lO0Xq4OKph0T8Fqn
OhODsQpNOR2ytgQpXFnR4W/dyDnFjbs7BdjOlmqYSyNR7ZZR90z5kiRSl7UCq8HlZUMPUmqfl8vv
Sm3qkrUQ9oPgBo6UOsO1PuD4Pp974e/HFuHgkfgF4o8Ck/cmaLNmBfx02EgbeDWvKbxn9HuKfgAN
dclqRZ+ZOgHUwcHmzIx5W0Jp9o2CTkYZZ0CZBiERZjaS/borePI2MoxSQepS0qZZdZP6tyP0oJj2
mc8IO8jC49qNUhKhnGZ3f6Ptm1mp6lithe2OdPr57WN2yAQAypocCylYgH2GK7EMxC5pZOI4TIst
XLujSafjTjTdVpKjv1IXbxG5ReKXf0DdmSSfxwYjaviSzzSfm+W99xm7hZO9v+Bo1wj0F1UVeNYJ
x8PpcJ0Lq6rr+FDT8o5n126073JnAr/oLeAlscRh8VZ3LX48a6gZqs0pfnWqMBg1GQ/9Odt/1M7w
aI7b/y2TjkGdt2S/D/eOq5yPUE00BC0BO7YcwQg4kQhoUqwH3WbLu5/gcvdsbSNr91k31bWZ1Vlf
CxLsu0GeaahZEQmTo1HOMdZNQdpEPJMQg+sxqD4ednxNcRwmQrv0klJ9OdwI+c59Em9FVoRl84ub
b8O+uVWfhYDBRrCoWJ+BG1QigVCGonp1VRFJwBH4omMcmsV5oL9zsv7EJYPn0DyMeygGljEIxAu/
3gFu4psVneAT0M4tDAuSeVUEamfVwCk2XzMDaqZWqJCUo2+fGMhQLLc8LnrMbppHfKMSpJ7OrNL0
GL12ENS06QhORSeq9z/0me4D1tyequN4IUzfjWa2BegO61X2BYRH8OPtELqg8jQK9KdkLc6LmMHj
P/rwS0DdtTy+JElxz43YI7OIXdGneZH5+gSF8L/MJaSJGHlCopuCW+cbRn083xNAdGwI5rutTPl1
67fCg8nmEGF2BKC+DN1r6Qw/R/QVJCOuCBt49CygAaDTiWAf4/NnHmo+jx++By63MC8/86JQaVox
Tlfevfr5sscN12kz2xrlqvEbMVbS3oQ8c2gX4ktjB0/PW0fsDajMivAHVRB+apzJ/77WtE6DuVXe
AspRMGj5FpbK0z3RFXXxTSWaYKSCbWXEbuDh2pvC0Kly7+o/8P8oMLKIrOurgcsHadfez+g7JxD9
8O0zFNj6RJ6rtYgufgroukd34S4rt8zAQ7p0PlP9mIUn6jd7pnQk4eFXnFsbffc2UYrHNcgqFa3F
XoBLheGMSlTVh+M/jrjciFSxcMRucRX3uPz/0oTTZyacQq+HNE5nbeCPYLRQHWZ7TlZIGIrxF0vq
7TkW7ErB98tjcVVwYHuRAMA39XtuRNl1TKOnki3LGrgitnwNGO0w45VfMe0p4uAfapqzoevZBMx0
MqktVMnikYejGyOM5hEqG8FT0704EH5YN2I/TcWV+h+bGbj6paZpokZJh+ov6DygTHKwxg1R7ENL
7on+rUNDkGg9mN9upZSqmh2gavtJmGVwH/XKYnZc4+Wnj9MT2M+gPRWRxd2O3C0HBJCgZ7ZeQz5o
FHp13gLMcmvRy/wLHLW0Cy5N6OCm/0xvE4XMuLhCKszsOu8lcbgBp/FQG+GtoemRypTibYGiMoNL
BiBBtekVlJs/XcfegCsKU7vRCudBfA6DtCqdD9nk7xYJfPR/I4ce2eUm0FSyvAgShwIFv774R3PK
JzKgPNGY2U27GCEG6doE3Qntxx09vmJrKJhsTn45DrEv4W6/FxJZl2tMPCloCMIuoWFQhn4lBMqG
oVZ4MJqwKo68YdiJYS7UuO6j8maNGagEACKS7qjRa7BOmpf1tGoDIynvdHJtw9ExdKOUpn8QsoGQ
f366rwvI2vK4xqjL+TUVge9EdF9nHrrxWcOfXAI4vTl377eCdPv5lAIGP5CHupUIUJ6fFwPtbV0G
MacY5XABGq7PyemQSB5j2C8g0kGcmvLr/fNrio176hsK3zUjypPJEOomPjvhulraS2KhMHjBBLnU
Z+Ebh5XMClb3H9/Grvc8RA7e3gFqhBDmU2KopcSk7RX9gFaVB+qYgcccFUFxymPYMOyf88s8HcnG
FAM97J6yYAdlBHTyhJVex3WeQ3r0o5tCOfu02HC/6iuaLUjiKiV03+AF6XvpOruYbH/feLCPXOlN
fg7oiCG3IxHTEtFW1L0dhv6JnBvQXmNJl6/nDrkDxFBPfegct/T0LZgj/uClr7kgUpLUlEA/LzVy
pgl70REdIYuh5cD4kEpuA+5XbDmjnubVQuwlT3xfeLL2nO0MRw/nbpV6sY2SiCJENp9xPdy8kTlT
qRrlDbf6LeLDHVf+BhkaJkAHezUZ7Ns2rd0efpnu71sKl48LA28lbooCZHwWYy9aD6M2GG6PQQOg
2Dwwg7HkDqLnRJdudawubwrNhP5aLSiY1yOmxqt/VB0NRjs1n1jZiXqsEXbrANFnLrrxnNY3toPr
H6x8nnAtqjZwahK9GBlIUDFgxvV4IQDemkPvE6NWawdvDQYquL/lLnCsOxqT3F+RBOZfnkGNYzsd
k53Nx3kTOxmdK1MVm+uqnu+uvT7UKK01fsIlKxEywzd2AayNZsmH2wq+xtVKLPHtTB9dEOQyLft/
pQQq59zufB+3R+B4IFFfQ1N/xJATakcm5lvzjwF3YaHdCLpx6tMup+QPtgWcKnPewKxjoQHpSCnL
RkZK9nY/83Jtj2AHGsCjnQSNaJI+ikBfJPILAzQevx2ajLO/aerdfnpj5NPlW6Nb03KFYxvUFJPV
WJ0Q124ofBWJ5U7pU85h9i1TVITzugMIsTgP1qNG5g8V7/sc+khFPTJh26KfqaUSNQ+JR/LmcFzm
eWCYrGhRKcwpto1l3/uEoHdpr3moiGV8EbySjzidjHvvHKyz6LPY3SOMZJoShoAQZAoeG6fbH1Af
8ZI38XgHLXSQF/TyUhC98F8k21KM+K+ucFLXlgH+QDUL2ytAxVFMSNrllSLv9XGCfQCS+YFwMEOn
DqepYyV5eEoRrqMaTMkSvspWWJEZ7bfFlItU08ntL27Wh5Biaq3+WXLApyb4f8SGKTFoiTtBXRhs
bW5mGKfP3n9y8vrRi2yYUqPdhUfVrMgCYmt0E+q75qeGHPAgJn7MsHdBUFC1/hN3jaCvDvgkWIUb
xWb+a8aYh6fPwEmCA/nzg2j1r9F84OLS9Yn0P7RzIK1IMoMLNf2mYK5D9jG0IdhYSgqEu/expBik
3uvrtWjJ/rAENmlj+u/GAO3eO5DbnpGSK8afeRXhLnbwme059vm1PfbTxkq3vpoTB03u/tidgHjh
cWA0mQM3A31LXjwR7xWuytYn6maRwo/Zt4wE+Z4WCfj1m0yzybFqwnq49ZkLw1NAFppA6tr9FdRO
l3iY++hulc6yS1xVBDDQgOOqvRqD234WahwVdEB8uuG2ESca7JcSl0OWSE27qMADIFyUOqse0l9X
+E0bpklVyzoWEyY1SOiF9ltab4bA3F7Rvgit0htzd5u4SyLgs7V+JPMJP/o/dqTznwsn8wfQrWux
Ztf/6AmvqDGyN9oIIKDHAenzYQXDpqlHCHzmxZX4DcOhtj2SfmDubmwufYm/cNDxLGYgB5W4JXVH
Hd5PsOgEgsBTts5+dVen0BBtTEdYskeUxPO3H5+IGj0pdOETlsNyccy1YTdCQbs/JyqZMMOsSOmQ
CU3Xm+PO2XwzU2qTt891ezs3/p2tdcNuVCEYSXnWnngIKCgtlFibhK69RhSG2W9TrTIMZ3wAkEnd
7eVNDn0C5wFj+cTjmeLvmURpiNAjWVlIke0TZ6YePLfcL6+OCfW2ViltMhqWzHqOuXoNiuCIGla2
3DOKfaULkyHXfg+m36u0G+ampEpuDs9ZTcDA/C8m8s+ndII2m1vTqzPpPEv1AzcgiEoX6tnvRojl
aEn5Js1uYrofqOiT6pe7aMoqQl88TZtwNkkmsZM446iAllyPukLnO2R56CLhbJGAHdjmFE10XaR1
jHD0i9FgnV4Dh7lQill3h43EvRRCPaOZtYObFbV8rDDxCBtrpLRj5gvJW76Ej62VziWFRm2v2W9J
h9LC7VUiGToAfUhVOzy0Ox7yjInysrynrFQpHkscx0ig+A2WgQEqkOOyTtoHG93WoCH8SShmtF49
szN5mApGewzIeanAgiCJ4K8OlYRR+bfr0YdbW+Eg143G4Kp+WTWLKgUVOBWOOyQQjQzHZMPafZja
qonONGWUJEmarlPyaZsBmlu3gOIYKqjn2ER/WCARTOKUnsIhua5EVW+1suCgwYsyOtiawd6C9UaR
O2i+2OmPHCcyw/f6mUn6iKz/ySxWT8rbIwtK36QXjrxZwptncb9GQul/cLsZLjd3WPr6NcWEs0Lo
JN5+xCuo3cY9VZZSJ7LAbah4VXqNYXGM2JiIyCeuD++xlFfTsYHQ3gnHn9b23WLLPBWj/i1mDN07
akLNPCTzKDc+oNCOMqOO5w8bJtOdwxsAoz7jev1vNhvEylH5l3MscGPoIsuBs++P+i8oDNTa16Kq
r+tyf/0/Z2OuqJsxcvozwPLt/7luWuxTIM6WHwBD7ZuTnOVAylUcC51ynWb43uXpOyWMtciozD1C
staN5YbPb0IIGFeveUd9+WZxqYL8UCW2brOaNTUNmBuE8AGEBV27DOUEdJ6lvz6q2XRif1TESO29
iYWtBrqT/AwibXZ+knfb0iMGLn/VGLu4d9RxS4icfZY6VEPi6go+eMelky34UY84JP4i9Tr8Un4e
a/HRU3e9l/rdNM0CdzhTdki09ix9b9iq8Hl20dxGJhqjvIcZ+NAUPGU+vZv3L40M8jQef4YQYt5i
G4dzvRftbLUYqujijCCjUSPSDKU5Kntfa+6YAhTwuzHke28763P6pd/cXkvrLvYYjEe+TIEJu/dW
OfW9wuRKc4QUIP/HFc4sPxFM+gqq/wz3Cha/mW7mYsL0OOf1gKSxpyxUSc+mzxv8SKpBWI/0kMlN
iY8OGcbRmFYZhFNJUA5Y7intOkUvxAdSxGfbT4RDDLQnXc6LXvj87JnHJLcdqxg9pi+LyueI4YNx
NYeDQ0jCgLwQ/5A2gvEImp4KtPZoxIK5cuZ08h88Tf+rhkh0u0tWlSdJDg1FBXuvrCL89wbkjDut
O8S9o4Eahn5rPkXkhIlPxATKs9Jk17MYDGfenw1SeuZC/QGxMCwrugzuLu6n2Ecq+KkU3SQ8ZCRS
jY1jaHoxnYYkNsAF4aAVa1dVqk7adZITjvIVGtfu3vqQIMVGPoFwnjtY1mxomlo4Q53NfHSLPSvS
RaUXHfztQT1HG+cB/y2DzB5ylk2oV3nxnXpnHazsPlKUgnR9v1ectGSc6rXFzSXbVv/nmrMULj7p
2392coRGkyWhOihf554VczK2kmRrRTPUeOqJObNn/s0nt5Fr/Ovt/uBQ8iX8ZYG9BWGXfM7v7ite
pQzvF8+xHH/DErCqSjLiXXhwLNbZvFtfxtBI3TTbyN4L7KbsOKpRyqrOxyTvTyY/n0ysLhuHCX/L
ncoVGJw7+LbnN/QfKosDZYw5MG4XPnP016BFv/yeZBgxDdTdeab2uywmokkp5TBytaXzbuT8zer6
OvTWSXHlAxRdNJDLZWlvkJ237xb575a6sIJekzc4pQLBT4htXXQbmC7LW/eLd/tRLuzLk1sMwpzI
kBRjmaO5Zoe5/OzN/ZL7M6HVr7T+uUTD/W0iKJwO4KvgUS9GzMcTzzmQ69BVU864iJfu3fBRpcVd
a3LNiHqOGrVaK22LK/3lDhQvb4rzUmop/VlEQKKT80JHiFtQpMrviHwNSFcMdGQ7oNbLqs9NItu/
+ZM8i746BceE3qteSd/ADCnRjc0Q8cgkU8v3brvarxk9l9kht0VLL74X7lmipCoVeki6+vofDlUf
pCUpPyMbTbWAVU14SfMdku7pJ9p3A3Wp153DCghWBWE+hygpd1Wa48NKrx8XMyWnyKOwfe4HtGkQ
L9hPy1Vc/UUKMNJk8znezzf7Waqf+rKAYrfJSIb5SbsToRxx6VswQ2d5/7v1mAfk5wiM6avYMFF3
In5cWv8ifda8ngnihOs6gUFPxWSjo7tvJCohy7JPckH4raLEVNwCjhruW9jllvdX1I2IMgQOSG8o
uGBgONYdP6K8vSrzBJrPtsnmBBE43TtO5eqZe6n9XZMJY3tg0kbN3NufvbGn0ssw/ufhobcQwSwC
Fr3CGCd+LsQkheVpOPqxcPCtSA+dUcQGsH9POZRnQy+Un+qZq2LeZEEDZQEMM8efvS+1nNP8aCD7
t8TPH81K4ac1GzXJwwvYrEoVj+q3f+j5/h5jPQbYevFk1L4w6D55JM4b4rAcquAOuJ02AFA7AFvj
upEXzUwMzetJkI77fd/ZR3PDjeiE7vITq2GgwLop4mWQufpHcQoXgllOT2uy+4M+/s7dBHydK0FM
/M1ysHZRP6o/ygcgdQdbqSq412DQ/+XD17BqA6ml514SXFtCiaZKgfvNKsiBGcr1MiJ14t5G1bQ5
SofR3dseJ/tjQhqXn9xgL+tnJrC+pgIDWVKhOMaWJvEc7VHk7f6Hhf8o2mNfyUVb30BBIcyUmvga
u3uGqYzzD9BmJY1qIBGgXQ8zEi1LhJIiU82leKsQqBfAFyBM2IFHU91rWzeOuU4MXjXcfOVmldsN
d5DmrWPypK4aeK6W5633Op6FcuMmJJFY8ZeNrXSNQXruOzx1Iqq7QViwj2BsvQJYKMR/A/976Bf7
s6p3vO9hir24v+lYIcbUtRwSWiXf/kvhckix47iwA0I+94aN4qW9oEKQK4l1qqm5auW7Mx+EtbTr
ee6vmSXkoOI0Xd9NW8v2yleAz0AInhLQiTHDw1lzMqTZ4j3OmTnzx1M1dPoSDlnJnokHpzGU60Vn
hqvgicmX8UiBj6VUquzk4EUZCv4vT8olmexIRETZGBW2TMKdkffjRQjg67ddNjJwL18CsXMlm99k
RhtIzOWtCe2h07/a7ThQhoQOkR9g3X+PWLsT7nImPHBeAuwXN0zsotDgZjodFx+wPfZYCGpgrwmw
LNRdqRROiXD+yeWo24guSAT5SKnDOjYIpsM3//nU20FSNDm5JxR9ZFIM0dBSQMBy6e/JlzgQJbFE
kBdB6nP2/WMqlUnBmx0P2WFRJRN5wOxuKjGaAVdJDtYQnzJali39ctowwquwNFhd+z1D19v7JCwA
U+pE8Z6Zib2H5l0ZbrjHbtBR476dcOg/OI5nyLzLziRRKvOls/pPBc6PxHsoCt0D7Fskv4P8N5dI
cdFGNeq1E4KNRkdMGOvXXsLREJPekIePX06ywCL7Q3i44pCcm+e5t/phnSFpbHBDCLv0KX58mZV8
VkMLuwJmgzOjsS6h8LvqUZi8GWtl/qwlL7AVr8LK1JOg7vP/5DfBkNnygoufnmJhv7W2WSApKTDQ
FzkIRfLk1tv7jJC9QsFfhylOpeRVpV4yfKcmyvMwJefwOgCaF0TTNAcgdiu9IPn/5U07osmS/Mjg
+f6nYVWh0BnCiAY3lknmaPAgyhhkW/L6jsZgx715UX3zh83EXSXKtkyZ7uybQLv0v+fkTfSsDewl
MuuyfrTL6NQNJYq9iWtx6UkSpKkKkTkreFiKeLGsQatf77Q8JVM+N3a46oUv6cQqjPPJeuOHbgFd
U3z6anCgBhvCGxUJTwhSu5xO1VvXTm5qnLv2sC5mNJaGYf+bepd2vxWHvwqxpqq++rK0dIOwEz0C
NdnmO5ZRfUB2n1RCk1V22JxuuQ85TfwE9q9UmJ5uAYXVFNgnA3umMkm6CZcvDSYZErxTC5mCQ884
c6m2uR2EKgb0Hh6ElSfRHZ18Q68qdoKJssYo2tNBdpIG5VlcX5Kb2jb8WrUqtXdcup4fH9RamHRw
7UIq2E7iXqD6eWGV7Rc6wKhNK0tqtuXFHFuf1QG6pTtfeJ7aBySO91VJ+fHutcJAlIYBL/CLHTgX
jXxg8JjUin0BSzcqBK5EVqUSMjvCgSKkxsbl18ET5mObvYcq/5e4DtX+qQlLH+XTwohZuX5+B5rb
RUDR+Wdb0yVoo9Ky4Zph5g+XKy3LZ9V8ZGP+Semj1QHq8qsUOkE9I6oVd5kCHuyibeaMGwj5Bqb+
mytFolYKrRUb5BSu/+TwM7BycePVO8HUzLHy23uNQvoq5Shy9MNgSCSseBmVgjuQPrNLbWA6Z6SL
I9XochJfwHkCPVBwZtCrvSvCnbZBH/9NfJx23puIIG6pcHqYDlhjvnZb+SJsJ3CCnhqh2s6X5AIV
XH190szpanERWBmUBkWq+5A49PNwHvFEy/SFPpGX4M8lFOIKZ/0kI/0SuOHKqEqQUaF0e/r/pCSM
A0BzxSFqlefXbwXaW0T9mvhIuo5vTeTCl3brdiZL4XY7btdMkDr6va3AkwOCrQLS5EYGFKBG8Em3
Ji+8IRybQv8RA5vjLRHyvf/IHG2mk3nKl7iXvzYrWEqvA4OPLYZyzIoOTMmKbwOaEjJ1tGoAfsgF
g7opgue6AwoWg+X6KpjQJ/3matB2XYFkdm/uMv0vDu9DXituHb4Pf1N9KIZeCv15g3sBkYiFgOs5
3x/AxsC1GqXlwVjCcAuRHwDAcUMW4Te+BBgxkj1/aWknMeIoXCb8ceRndF3MuME0ZZ2TmQI4JHqn
P6MPBmGK+yEhraN7oV5wd5sf+wh1ZJVE4fz35uSmTVMkMssjeDvZSuyjmeFXCd8ehl5EmvLcZhJs
6lgGCuX/DO6X2eYuqc85AebL+3vmwi535tmgxjjTq35VAyrulpqlnTcesV5Ap4o/FjakR7yGvsuR
PNXGT6AEvCaCtcCDU/aVmkgUYldeWBvLncNUy3J9TwKONETnehfn0Secplv+j3ZlkLFNWgfojruo
/DAObvjU8iJuSEc1oFnMcJC+OzyYC8jc6S5pYaVa8w+tYOeHnMsrNZHsO2qRazng+kMbA4UOP7oq
Zip19IJN5hRHXINXCnlxTwrucn7qkzskK66iZ1HBRpeuU+bV+QY1Fbr2kj+xGPl13+KvyXIGIWy3
pDpF9A3+mchwmK+eoaEw+u4iUI9u5L5kZdResdbHfPG8naZJhKfLozrmrkqtOtUUNGF7T7z0JdAr
kDha44HxVFTXYAMtVBVjIp3cxVYnXNBCnbUNhRTUysXZ2zcolivXabreIR43P/QzVKUgsqTgYrYl
I7diR3O5e3VF63iEgvB9IBnpngsDx/a/MTNHvsd1IvjgOZfIquSk3AzefNQeMB2NxhvHgEiXIv7d
ZRMiahvltuJPy9Ws+SttNWVYBzJN0gwXTyeVRrJtcVtRDicNRTJNHxkNN+1BVHZMWBEBCJSLapL/
AlN9QbgzlPfn2Z5KiRWN4TWppMQppgJaTCGcmS/IRGZRZnbsp6R41epyLNChyPSe+Ki6VQ5rcTJU
1xU4sGkWUcqPx9znBhwCDREp7s9eOkBiK1pE/XgtOndS1JeCZOvd7EyWu/fNlyvACY5o6/ePDtGU
WKZFt4wlMUu9gmLyLMV4eh+3vT84k+NNkmWFK08KRXxcnszOmTygi0SRAtkOy76Bdn9tzli4fMXX
wv1uMs5kMXW2sLiUyPMs5VS4vT2gR1Bvbt9945OMXABQ589RBcA3LwtpT0OElL/5jPFvDx3sC30v
0EPd54x5oe7tGdrqo40B6NgIv9kE9LgF41CrFWZNMItvkOhkSlm2QZFISvD5r8WeP4YEFaal+ynM
FweOm1IByYO9ka7LzU+nBLy+GWPWVLQYWUlIOcR+5auZ7iXyBmueshgWCcZJJL7uDqHLWmq0HsRA
cueAC7Q35Xa5JHHZ63YAGSQRQAq+OgFLFofu1YzZuAqhZOkmlAXzzyLWY22aZapf0nMdedMDTAWz
PvbjtljGBjgTq1aqImWUiuwn4HkBE9nvBg5jclipF5IE1a7S0snYJG840fRhRRkyWGtqVOAjR9o2
RHHtAXtrVgVs7hL5zQRC9hp7rx8RLNuoSAtQVV1djQ62XRXbUq7mStBr+bDJ5S87pVqm+9xfpFm+
7Q6MqhU5fTC9p4GfAJ3FA79SL/cDaBXfX8Mnaq//YwzxTUnfivCNM6SWfKHn6sitKwtIzcZU4XQD
qFkZdumpsKABDAJSQlUwUkPRCzyYeNfx5qpWS1vM1StGv8sfoL6aqIibuVn0TMbsBMkC8hs2pmPO
GACCLWeal/sLTqT4NPVKXd2l8TQ1M9jgyZaBQyfPrpMOXSmfa7akr7MN5MbmslXaJMRqC9F1B5K5
3+uwpEzG3uvdlbvbE0wMnNS2LYQ0bmbyaOvBPdxXav1oWOloy1qNSx36HoiljWV3s3PhlY68fp3C
lq1y2gceABnzDa0DdbfQxBx5kTpR7k2I/48RMVjUBdbaXkg4d6VDHfBIxkQm4wObFJDTYVlAa5oW
se/jsNM24KDLAvzxJA6A0dbQDNwfgwUHwrZ3XiwC353H5ISIOfAImMtFmkgOWqTjwcdgkcm07/aF
HyZA5wzo1eaX2m/pIE0CqQFdWgQwI+wl+pJy48PC2jqNUDn7n9XMc4HYCnlB8WTnqECMkV4VgteH
15raaPm+nkv34ayONw10lJuTFH50yILyWzaciWgYVA6d02f7t8RQgyJqaBiB0peJ3QdDvSz53ble
EZn2QwIKbJVe+oBfRsVxJDnXny4/6YjeWKJwPSgahkQ9fahrkXCnsscXZv3CYuMXiyihhblDjR1v
vxonT9BwBgw9BsX2UcJQsggtnw0p09QWSCMErUpubDsrL/H/9GV+FkawaHL+gNwJiJawuQTGVotw
PShxBfgGOFBMebzrH3cLvspbxePby1Ca4zWSvZiCVkEMfHrCI7LiZs59TmuNGWvDDmmUmqOEtVSl
cQgTQE0gauz4vUMU2guK/MxIQmi+TT3ZgtH613jE9pwQS0PvETgEjKOrwh4W9mnTJW4Ug/Q5Pi4u
aviWNA9lttOM0lwRZedqW9cZaW5ZOz1llLxE6L5NhSbXtA7LcCDS81FP3qusbpiNf6Dhj19stb7p
dQDllrZVw6n5XHMPRX3u5zCleXzkBroAXz3ErHqqGiiQx2oK8ZAWD0xbtd5DdfkvPfbRfRxSjZ4b
AYMQIqQz7CeX2B9EioJgxOvup2HpP7voPOJjbc4vA9kXi7+vpikfPULIG8HnriI2FUU45hx/7wRQ
uXiuA6KqhrWmLU1lTBUPFwX04L88Fol9UyyMgtL1ZPvat8MpHDM5cdhcYPeYYtU/6dTxGVt/4Bo9
1m/HaYouhPOyCNhy5Be2nC9a3Xuhfsm1cGDlxz2ahYrTh3CXEBZGU1fVHKx0ULkOl/1YbPVOxhCY
n2Hsc2Rmp29O9iCA7/EJO2flW0tB49XBadpz4XCtZYPPHoPGIWH0oCtygNfDVV3mBxBXOcCqQoHj
o8EcLilqQsWUm/h4+zUU67WCGfdsVrZIULPk5uT5hjnevsn9GD+sS3cqxuzN/8RHB53HiMyqdpZ+
Vmo3VWUtbIap5PXdP1yx6huiGGSJTWFwUppzUM/CmFeVi2TNC3IyeFbuJkL8Ow1UK+rFV6nR5+xt
PBZPlIW9Jm1dek7xlw/RATRHC8Hj+kzR550FlzkookO4KWYCQ16iDEnqbBtZWzn2Ye4kxJnrF1Lk
GeUYHi/Rqc+gZ4HeXP4UqP+bwja3ebt33iVcX8UaGwsJgl9BrjkqdJ7H04g9sD1rLkYsEJ/lO3yE
kcfchUU/nxRgM3MPr/r1SkrR6PayQ4x3hSdMLMM8g8HeiAlMYkHYAZtMnVRYrEcfFvqRw4ei7Uht
Wb6WkVK8V74KY+0hwGB8f8mb6KKSg5VGxK5IK0BwEm8GwS/2LUUf+V6KQ0Nn0Tr1x9j7OgBhHD4X
YCBP35L4btY+C3u7AGcGx9clmDOmnvUYDoHahSxcDbQi1ATyAnAOO49gkMM2Big0KRXthVE6CUz1
hPwwWQUUW1QvIaRVBevE29wD76Z3WP0WBHpabZBMxKVHV/9hhGGZa0lBByvAru+xk0HyB8M0/bMt
0fOuPNTdYPg3B5k7wf6NsJL/17BcXP1/qwXt0JWuIPK0r5C/OqRi38zx1x5ApL5R9zhVx2CqagB7
WxbO3s55SJQRBTdZh7Ym5lbb6Jv1qkUHuc9kXRypLEtB/JDsH9H8oLrjUcJKjiKeMljWqKIW9ERi
iTYpN2jhm7mj2QfxdCaO656XuiEJjhkQIGWAYj0ZRaG+dU9ArFB/8SrWIa8WKVCPRFXyt24AMBW3
U5+R4JaWeiRO/FyBE1TnJtV6oHjgSrUOBbHtFGQLpbn2VSjAj20lqGEsaz6cA/i75btbeGBBuy1g
gx9l4jPz6vEfeYpKxQsCYX4JYgMLaFrX+Rbom6z5RQzjtEJF1+isLABLcEcoFI49rREwxGfMdDMR
zWOBkyiiYU1+bmoQqsujGt685eh66NbE03Fui2ESMjrAgndCphOdxNixmszMX7VRXe6UwW5T+jpN
kFSBzcC/qZSyYGecEEIRrVazz6F6m4HMu1MTP00XPEGraqCdnoT/XNaxGUhFHoZkpB6XKzJMKdoi
Mj4g65yFINl45cGTOUTRyo1ez0OHLZ0+TKZOWYvd1AXCX5bmEogH5cxvuxJkV1JF68ozOtJ+q4ad
dzaufPLhoe5tryPAm2iVv2rguWEkAaqnKNgowusBw4Pqk/oJhtSva1IMqeKYugBBOF2svnuuTSbQ
HKhHQ/IZXf3Wx6mzf1HCe09HOmzpmNZjE5ilullBb1LuWV8kIg20NnddTCOVor02Yc/ADSO/sMw2
YCTcvXinMWJn+naue9fvGqRYHv+q947uUuSOd1nesuqg2jx1mfCiv0LC9eymmXGx+SrKAqurYjUe
nDxzFuZsO7U+jBe5pJPsxerbj0A2V1usSzuMwH8eBmfYEmrrHepot80LjWQUbBTwYwtUwFyWtyU1
MB50nrmHnYVoRa2CFoDgo2GRiSwooFk3XYRHRykA5Ycb1O+7zyWACeGQOgSAiiGUl60FAiMZwspz
II9Jms++pPyxL1/3f4Q/Z5IGk5/6aEw403xPIb/xlvzrJJs8f74s79L1w06tYQIro2826ZvP+q8j
TTTm8Dj3lUzjrrQ/HAPCiE/I0ejby5OHRn07h/0xOLGFJtR4Zlz0tjjAIbz4cGljgC7Zvdy8g8zx
dxBvuuW2YRhmvWkISwXeeGCg15e4d0gljCqeQvUkgrZb4vw2otQb8hI4tf0K/oIGZB/fEY8wmtYb
A5EChi7PAZDeZHY951Ac9Q7F6QodOw0PfOS05SzCJzOdD1IbKuRAVtwUK9+Wzj3VmtPaJObgW7QO
NNeRPc391BPYzbGGBShxjQDEWrYNRDw0gX8VTjqoDDNxve/Ash+X9kjYN0kS8r8iLHwdlRgF/vku
TBJUtTjnVOg8rhqaNUCNBebjLTX1kTDEK3/Irsmyh3ipE+evwsLX901AW6TXOrsMWmLnOeHgbqNI
gXzMDg1esi7FpnKZr3xOG54A9oKpqOHUrRpGPXVy9n793HO7RfSfv08s+0PKrDvrajkYgJ/y2A8f
tbMneiZiAn8YnGxR6oWkA04RJAbNNY2pdD4gFDvfMbawTVFBaf++U6pxlDYkWemIP6ECC/0QiUsg
ogIe/sckIHo5W90qS2O2VHGW+KhycaNNBbewHSpyBy2H4SBlxgG5+RqnmDdrUKhgZAS5Te12J10D
frNJ8yH063ALx8mEVUuvexRxyRfQtTq7LrOKf1XhB6GI3sLk8xwKnVSxNfWP+VV974bveD4KUWPM
HIMGeuzuDG5YKVHXDGOpdptM0h4TZNFrx1zwXRGmTAe987YFheqrtQXSDeHXRGpD9LJQfCQpQx84
7+XJVZt50fHl9whsi+a3GFK+FFY62ymtpyrFglPSlIEJ6gc2Cr7kpvjjTabJg3OXayMFK2qF5El5
lPx2vGzDt31yAQnJUKilX5pY6gCfAeDcWHmHWCVPQDYxU+jU+yL6N21v1ZR4Esrqxe+3LAeFnSix
s96lxcrixk0suoWrgLDauDU5vTke7POCqLqhEBGSWBgOWOnyxlVbtDvaMx2k1Hl9Er1H+syVlaMG
Xl0OWO1uxPoJDjApoyYm9CKT/daSvvwmpw8FOWMb/v6zI8FcLXClu72wexGUOH/i13mDc4DmO2zs
WQFJWOhAGY7fMN0X3ezQMh3SiO7TbSiApPAsdtmI4OITDQEdLMfuwblL/lSbLZ3xaOzByKS1XNDx
Km40cPwMwnnS5u3Y0BglB+Kntd/DhYibCnPqmnKl7puw/C8LpV8vzpOL54MNt1aMQL7eHxV8b5Pu
k4k9lrnV6g9MziEF6v2WCwZut4gULTm6Ncn46AEnE9Xx1WpUJ9xpl9KuQg9CsjewlKX8m4moth02
iMwbfzNNgvIBUh9B4lYd/cnxHV3/RRb+m7uLbFnamfVKc9k4AOIQRV+Qo6L8CLECAxmstxvbJNKQ
hT0BIGGSu598vjRoX9JZJF/Q3wYmxm6jtyoRSHEo7PcWxcmcjKew8AqdminCzB3gTrhG9ox67ul9
rP8tztnm8pt1DDV0nl4dX5fKlzIinCP4Wo2O9ubwqB0o0yxp4Zml7mc5dSlyJDaCIem/totcdWAG
okr4Xr11ZGQGNW1Lw4jPju3Vh3UVBlcprFGYthsdu3n7npMvAjhK+yqYQ0kvRaB7pnjisjC19GbK
imabUxqG9If7bTp0KAd1Ecr2Igw8rG6TRAizOvOibhH2lTK2Wwi106IlaJylqmFX0knjWJXStB4z
7KUgFJPrM/jTAQUyxKajXf7vYY+ddV6PlIZ/Lxs+fjbgi93o+cnNgW0cph5vE6ZSy+X4X23wjh6S
DwvwKU4gkWthn9TK04K8IAEa7HOjh9L3Zkq9eFW+1Qi9CAJdoRgPfCN4GqFQcJ+61FJNU+pQJXMP
WL2yfiY4JOrHlY6EpGSsYGYveIMoeyQcbyFqojNABItoph3Ky61pwKV7L1NmyWN8HBMgC43h+s65
ayR0BoYvDsW7lD7Z/vKiePXzZNnNS1/QeyK5azc8qf1ve0fmTFwy464zgHIGR5jnUa6IBnT8TYaM
73VtT/bKr9je8Cv5mPe+i0Gv0wWBPJx/g/Tbyp3cunQH6E9UBoa1t3awe6bwht70te13L3SN5PJl
OR8yvo3vzUUJpGbcr2SOsHmRsKTxwLrylJtghINnzi//6NRcoVfSHKeB0ZgMHSygW4kdCAuC20Fa
djBlDvaui4MTtkXX0oeYXM4mc9zkHxXrsj51+p/sNtWRX7UyAANy8RzF0C8qdBWk8GJbXZN9Yx4y
VojmGBOmLrW8j+Z2wurKRnvXlomCC/15eYY/E5g74ts4rXQdxG/RkCfLk+LanfiU15aMSZzTEpaa
QpVo+gqu9rfw9CwGH+M/jFDGVBpgDD26I/+lHl7IpYbTIJr7A2Wwcx6xDcRwilCc7+u0Nv2DhlFw
7WAtLVRT3W/lH97xZ0h0aVT7efzdMJS9LH1WjaU6aEHVJx8B/3yq1Ry5lJbOfoJ1rg510aYsTCTN
oppzcCvx97LB03HygNRMhVwDGqO+GETUn7oj1iRlcH9tOr2Nc0gCuP9qxeBMYpCzWwRf6k8EqMIA
bwPbOFp5ttLBpACC0xkjmJxtsSOVSvoapVMiKTz/u5zX54kB2/dgf8rz+YjwRtMdUMTF+U6Te34p
5rBZOoOW9KOD741Cr7DQqS4lNXumYnSm1I0XrScfxFvjb7gVK0ArvFPeNoqRPRlsG1DZSqZEbSkV
Y0iIdkV01Sr2Cta0SIiOuzc1Efhf9tflqFRvlUO832bea/iMU5jybSqtKCPjIbiA0ya3txpQnROq
HAIdjmtVswUBYkZvjsCYlG9D9fJZYhvtGoqgioDOgUpVRzSJDdsQm0OiZZPPCnGLG4D4htP59uMe
LkijSFM8IfJvAf17kSI55HtHKFtS0ix2ausgwuPIWygDY7H0g0kxlTniI5S7fPe2P8mxc165G7kB
L5v5g7Xk7cFP5HmhPjMXNIq8d0bl/CwOYGaFDfNDjXwO+k5g1j4p4K6QuBjTJ98vSTL3ArbjW730
N/y+UsnfaJDqQ1CYFfSMUMttWbaZV/lf+c2szuMY5XWw6md8sokS30PCotreFSCgarzzD2DBqlOY
sMrTzBJHSbCx72CkB242uPJcrETZ6dKieQ+IVFG5C+PBFz2Deitk2H9MLNghVE/kclEsEp1fhTN+
yu+wlStJhod7N8nmQNDjtc69zRu5MjBOL0AmhHHF48NRn5WnZ6mQaV7AaNqtAzo2MP/2DjvQuU2K
8Vh2lLa2LmOdMNMun+VP9E2ngnXiSfd9YYMXqJGM5HigIyvKAFnWL/eL3ie0AFwr1v5DVYEMfI8Y
oPHWmXf0Jy1VpsWEYcZUexM5/iTARhIesF9nOgTs5el6z/Nle+QdfdXpIyiSattrb12Mv/HAROzK
LzTMTY/SYjSOxaFMyS99aErbrTPR7nSW95MktRK3OZOfFMwMIpgJUlDf6Yzffo73zV1H6xIYX9l1
+DIYPZnANZxy/U4WQ23MzNfYbP/sQyelVNqZVZ1hh9evScwcsaToUABZAy1HGmWi6VrNMR4In9mr
FSLERIfeDF7NPGigPZsUkKk42xFR0P4gQeHdUUIjCCPoULi6bvhabHfq1EzDjvKthtGl+DopKyv1
8JimtX1rmenircsNFzg7Ng94sDUCXaaxqoPzUoL3d2Ad8E2F7WYKSM2ycraWF2PF540ISXJlYyGZ
zjDZijnMwX8tPuopu6GDFnF3dkU6zquaGFgaRNNzj64uEdWX2g9K42tQ7rSpBnmtPpeulXeo8yTv
HSKinUF6CZUY4x4uDJpULcmxDMhqX1bMAaN3gX0nny+M6warPmUDi+g5eVkiYYgsmDrl0EVRsYkl
DGqmpcBA4E/m5GGUOxbRGgKSeAtclQDUSHHH8J0eu+NfBpAIF3UW0zhCZnu5HNj4wq1PrgefrIoo
jd8QqudCC8ZOEG98Y302uabWarQQQpw/M/wkJVSnE2REyqMcQaDWteIoMyTdrOYPRaGo0FvUit7W
QaEQ3XJYpnVZvpoQzzyGpQ+M8gxqIXbim8lICWUgIaiLx8Nv08TEftyIJR/4GllkkRig6Cn3W54q
CMkGNt0C95WmDvmaZItK/TuvpEFN6Pw6UcPeIneMeWFN3oN8r+SwKYS2nyOLT7XbtUDoJgxJYORO
Q3dZbV1BGS0X4EX+I+dlvAOIIkjXx5QWrzTZkMwFODdcrRzhHl3o1Q7Vfcu9GgVMyAn72fxWDk3d
WQhWtYTZVMfqeTrm5UnVZBMysXQB/0hE4tV+nbokAYI1B5iao4Cp4NSn/hVtRYGq6DrhuBNYIHO4
ibC1xmfv/SAKVdtNyax3M8fYbOegVpm1/+UL2AZLgoLHwl8uEWJYTDZJddQL4un7l/QkKdp9kQx+
+LwQKNHj5Yapk9S1Yeun4cZBVKyzGPqPeZDNGrd6cbeMX6ZQXmX+ICV/p7ugaifI06+ElVDSOGJo
7HqRo7C1zeUuFTEE9mInj066GPc0jlg0j/K8k7ObrPztkdX7PFpYANlN6EQOEtAR+rp/4tqP8gi8
EYgKHbh2V1KmHEG2WIjlhfv6yxm6EwGqEkddi8KF1AFtGyQC43NEympYOC98T01G6PcnTSshlRDV
+G/1dLM1XnepPw0DALTUqB0TUNZtMcpop9q9OQfB9VQ4Odm1vs9fVKUu+Ix+d9LbRcqhGF5eZWu1
xtpRT7y06nOJ/rYM2GexCjiyADgt8lKkbtOOczC+xAMd6BRjrbWzQTxLPxS3FNUe50asGkyQZ4TE
fcHCFwCW/oI0EmZfdLVRQGB2RZnHJC+gETHanOO7L85eaazTiPSXVftHedq2jx1DWrbPB0OLoX6m
7XWmlkqWD2ialPu0oyYXP6JcAhWg/ofRvhVwUgji7NmoR3ynVKtjB5ZM9Y6v8RJy9mMkwvY12MNd
q6IdLTXyw5RGhnxOrESoNzQc4tgpNc0jN2XK2QKHpy7LIQwh0UHJhCcWkas3IrPaXYrECAKHgbTh
niknfGQEKovrW6st0V1V9E6mBeneXTBIAij1zIMqRStmlKm8FlMz4mm6GUFhkpysTKrKMSsGYToc
3sP5M/BaZuX+HtSUQKovVMQtJXuTqzabLrV6949F+zNCoQ3kZxXrFIe0X68a1WHmm8zGgAkN3D9p
lrrp+AtJaNX+hLsGXJ/2XA0Rtb7xAnETn4bE2RiJflwbo38eKwuM5YbqK1QWIMd5EGFRyPLJrfG9
dVpv5fHmOdp+XFWu2/FEpn59PRczMr8bCjQdHrlGsnMAFHwCfTH/ji8Ejja3y89aubvEuxt7mgvL
m5w4svN1I5ER/HRHCVklywFJZEcGfX1YiWy4Rjel+L2HN5nDcRcKWT9aNnjfauyPdB86KJDvkeMD
tXU0Xq2mOBW6wO8/D6WvB6A5dVzGI09GPIrNp6NRa0AuStG/YI5VykTdKnw6lZ8wtAZ7Tnmlk8cE
zI3fuh0jHOTFibY0V9hDo73E2su09Bxmrrn/X3AOgUl1Z6H9nlwLBXbHrOp7vs3253fF5aKDuFik
utAZ91u6m45tbNHusUGbPmrA1dn3xvxNLOKdsNYoIQjsyKRiug+WG7CqmO8mb+2o3pzTuyv+YyEy
J7+XLjSzeB9kOz9lMKcQPRSv6/L8w9/iKWr2ywJCgGsUldwdORD7Lphig7tWey+xkEhFciCuxttz
ktHKtxmUHFrXAguTv3AkOapyOC1n6HCb3vFQS0nIPYEyk/rC6HqRcLiudmItnjOONxsoNhaAN0Z4
g3CYBZPpquJMA/W1WbH12bfmcs93uJ+3//TEAYflTDdkgc7p0XnEAQ2dpETJ7/ph8QOGSbQ4At8v
PTzLJdov5jYFmSFHLIKKagkDuGJB095zFoGC6Mu8rePN4zCByFKyImwas3+Xkc8LTnWIQ9Uo3kwG
3R8IHj0MlKGGU/HglU7+1kkD2D3wOsHosaPuB1vjKBQWtmp35mPyZRkHbYwsxnZQ/f3nbk5hlE5I
6zzHEx/1NymT2j7uRbD3bJvqa/vn4aNlVfnVbd11wmV5OOgg2R3swSvyo3S1mVi0cBbyaV9KZKaz
hDOuf2tp8uh2ilR2CojHLQCbbh3B0X+FuLDrGw4n2hSYZ6eNl9S2Xr/n2XCeIckeJEQ+bn5DYZre
AKs6Ai4RxB1/cxDIbux3ibl4xLKPvK2fhzOovjiNEh3KlLiDEfLuV7VucIdjvaDOHWZkLuf3YXZc
16nvKCvAOqSd/KCLs2Af1UPspDdGncZNozHYQD7oI9dKKLGL4BQcmBQuNABB0QsOEOSjktLPX0OM
saDQ5tbvi2Z6eTyRnqdH2sFSdPNs49dSm0LOlV4bOf+KWgPpPUumY/aQEN/Xuc+mfFN44DFZu23u
J1G0giNdbIcOWQ6BRzTprQOicnrLwJVBZAl9QnrD+xh32A3bNWtVl4rq+TNPEMEjXe73DG/xxCPg
nqIQVjdlCplGidrB72KsrTmOaU9H3zFBAcNNfssAMKLBWg6kSx7AT1Ydt1kOlGJn9QcFfn8wOeEv
5Uv3hmORons9STysYa0HoZtEpe9PkB2D2CLA6/rFnh1OastR5SwV3L/pX+i4aagnUOFiW+PEEt4Y
fDYWj13HpoVXrlnPO/gMzqhyeEgx0eoa5pzIG2qYTzXn8zLVS1BiMcgYGehBbQg3vHbViri9R440
mkUSUxdg8s4nqMsdrusOr8hJRBvDyqW6E1h8gjjUWOZP49slHEUvAHQev+J/GnpXME0RsgQ/JF/9
CVvhvOb4TZvDKrRoonHFKGSO+mXnw6qZfssIBLhWU7fO0pQLGKGwq/+OSSrMGlc27//IvEXIY8HN
ERduBGrHKg+hMCZa/5eiz0/jnd9wYMdyq4wzU08poWrcJlqsVxD56I5e8ZcDIboF+7SpSTWquVCN
He4fD+C161ylSSR8VKDg5sj5ooUQwMhYuGLagG0yUmvc62BiyhDMo0/F1Lzd2fZuzr9J1zyOMbjF
mQsr4wxxxwKuDwXfNYjZYKrfWtoA0BnsZZddJJrEzEDzNVVeZ9KRFv0zEXrquOb/zcg1QAWQZU2X
WGMMNHZgLeZH8CiyEvsg7G8KRZ+YiiveIqpHN0IJF3NmfPDitWYQ6aMyKV2nyBiBdyQJ3NFP6K0a
3/bO1U3icR6HAEgsaPxzZYfcLpy4OpjL7wFaq0apKbjBWr9cx2JvguOKt1rTCdoOy1PjsVieyhX/
7euUeAeDl6M2cfQ0dGaOnJlcHe3RL+Y1YwukxGpyUb6Mo9zFALnvAjFAtwWz5tHldDON7M4knpqu
KHg2/hBEomqABxwQrlG9DwQOG5LcqyjjF+w9li5mxl7IYiYMSzysvFVa3kpZs7dwzhrfmRadRlhw
t/vl4g/YMBdSXMIEklZ0b4ttVPs63mbEhQB/IItuO3bQscrLwKcX20kGC1mR8hav8rByHQ1HKRIg
k2WiIeyp5lk1zKgKDrhEzrdRX1bM1CGh/26Y/S1iiZdUj0FGb15/Bui/nesIyUXDb+n43B95P5Ec
tQX2k7FHq78lm1Sj9544h1B/osFMGsdbuW/HmByrHdLBrWEpDPNekFbBphuEIU0p0Au9SdDt3VxJ
NwpRUtFBfBkTPM2XdqQQpPmopa92T1bsBFwLkdttqhldvTopCSDs4hWtkGy/Im15fUGLGaVm37RE
crPE879gW443cgJcgqOnG3TyKjQmEzN6V9SiybM1fXzSuC4AuL0jqmKC6e/miUeXwbvtNtcUay5O
1oC2B3Q3y3WG9su1pwO/o1mC2cKPgwbslGZHXkW2o6GoEh4wl4eURiEAbKY29FjrP27QNDVqlWcv
Dcc9w4MEsY2G7ZrUKX3qNEQX8X8PXji1yH8M2mZ4qIPDzVUUzftoj0kCqiX4zLJdACEWpx8R/P+v
fizgY8kt/NbL/9A3bKoosYDa2+l/HeJMYmRMUe+EOCVGChMfQ15tHLsUvojD7GcHFDFaJhBMtfcf
qOSFUzLgshRG2B8k96LevhZGGQCl4gzIjYkYxQOfyln0caYSJ6+meQ4/sI/fa/EtREiLBJF6GMzW
BEyXMm52TCMBq3MEnm1Rvn1Ubx0Da6wtC8ByRKRyKm6e8zU3TNLVZBa6oQdQPE+SrO336el7COoN
ia2PDTx8N7czxXDcq3ZklyfLGDkMLw3dcXph6uLBXwJfEtyd/X49f6WLMfl5dmp8GewLUPPYDWzW
EcBSUmanbpMCuPgXEn1TXMNKqjHVuS/6/ZYsM3P1GiQBPnvLfOhs4vlUIe6pDqbZGqmUzdcVoEqC
2W+s5vWr9wdhsXSnE1ZSwqh19KIIp/Amezns7dXO1zUOaGWLUgEqZyEoNUg4v20n/FxUEQ1Ml3QQ
DTF0DJIuDXDNAXJCru8q9pJ2Npf9+HIGQe2D1etVlozoZYuJLdjKhy/f3YxkT1XQyr1Ka+PEFXIe
40b2z7vZFClKhPogXhQmazodMbKwbsqqIPcUi4Tar/dlhVRakviaw1U8DckCG5hN8LrN8t456Fc2
fWOcmU6+NJmUHbxhuhqXcBcxwdROe3Y4bP05LFv+MyniQE4R7NVoOqciJ/u9WGwsju7csVpJZnLt
l55phQiJ9OXP/Ii/9NP3W22C5vHsIvvELII1E+Qkj4iiQDkM022+UMkJgiFQsyMAlnSdBrorwZip
DnrQGV0Y7/naI3fE/4+oJ5janVsEJnEnbu5gbNBvPkzD26j6qzkrNnag/e7dUUv1K4VzaMo38j87
33iYT0QFvn+A5gPrdGiw75yyJPHH6Vpj0nHYCcoCtikNTxe2Rnfd2pWvTtQ89j9i71FxcRvdfrUq
rUi1AHLuUulFJ1qoeWu2ofUzXA3sz4NeQghidbp0xRfXePgCm9nEZrHEoUiJPoCEX21SG1k6+lsG
EZrBvOAweR18Z2cUmLsqTA5vZFj+zkP5GA/V4HCiQ0iWU0F2/sUOcohgaJN2WlsXByEOHyLtQTNC
rIVzdC3bGNvTOUMdwc0AH8zv39fdOxP4NIDND25aTtWOPjU8cOtk/wHnjcFtBPDlMJXFQAUkfS7V
4ndKXGzJnx9jT84pTt+xOYNpttFgUvKHL3pr9tbxsNWR/XworbX8eafJSKzDNbJX5EHxhU7ExUkB
gR5bvUbVLyBGe0H40Rw0ffA/fZEqiRFksME16NMsw8PXNe6jM4F8vfdzufY1GsmhTHVyurodZOWn
fxNx9W5gHqgX2fSJQXnXj9IJffo3Qm5o1xvsN6Pt+bvhk+F4/MqDySfNTR0KfqCq0CKIfoucqncp
TfMCzTMXLAwrU6kUf09m3+AdjfpUm7G6CzmrLLmL4aEu0TurLx/qvmNRi9QkSXHO7owBbDt4wVbd
wmb3URAk+h5KLEKsFXFPgH66u1O8CG8xzhckz96s5ZduBJYrmW2LCw+KuQPRh7HsbSYniyXpPkuB
S4Cou7lpsXnUzu1oUoBmuPVBMBYqW93hoIJGjHaU0yeq7Y9Drycf1REePgS/S7JJa2Y7cF+bHW1q
F04eNw1xnMqbVrSadUPq4ePYNkRh/XOhgAC2Ch0p3iDYSGYGoBvDwr6vG9NDJWaeY6Qy5rMLf+a4
zCSZD/scdNt80wP8/ANJdVbQjiDDbNKKECFyE09GWuBhMjkKojy1/gZAOAD6yyb0ZdXFOBFBUBzV
1lD/UhrtIHMbbkA2iF1cGLIhZqYYSdzTXDiIPipbdzV60BxEo0cmIAKFMI5ANFb7qhN7RKckbhhy
xnITIPoLcnv1lxnidaeOtB7d2C7C4wwiq+r1mxX+YtaWV1/dWDSXWnF5C82ST/KKJYMU93xh3eWv
THTy3+Ok110TSsXz76flfMw90K90AXSkK5IIxfBmW1pgcPQU/n1Ae9/mhKFQkjebRJMK7Hsg1/0C
ed20VOiDse2AdXfCGy+3vscqV4g4IFf5cu/METsoV217mpNYXiKzotOPRzvTOhaI5oNWiIIJTwvr
zly4xCws2ciLLxDH88C6evO8+xY1s1goNk+JxYjFToJYEK8xc9FrZMq9T8cHHgtbZ2xXGp3q1fmI
QLm6G7kJMcF7U+0PWz8nAwsGP9d2U/yaPQDhakbRKPUgYCa8M0oUH7NeqAy6iqT+Qmrpknc6bgG4
wJc50RbMbfJTIPi6iCmOkfh6P9sGTDsMv4QHAJkg5OInzd4IBAH2QlMK2jdlJVuYyU5o4QJrr44c
Uo0SiUlCxpiaCemA1u8Pmbx1rIP1va50fBhpkg5ws8FbaTpASmT61lsHG69ulk02Ie+60OdzgSZB
XLJPqWrMf8KTZv/jv7XIJ7wQzWNzpPlGXNaLwgoyH1a/ik5XuX+2FF1D5CBpNXHLA7UujpWbrtbT
naNB69Bdo0EgSx9sG0tNNMBTJ2xrPQNvWmPxqrija7vfDI5Lm8dGG9EtU9RQ002+unuxWhyawGF2
x5ELR/0uWQH4QRBibLaVf4+nWzDWHpDlhz+rD6t+bSsAB0VRNbQQMai68cMQ+FUHTPlZQgVhzT2p
W09J1V/dQoEBC56buXeeXXDFk+kZWRUm1C0P9+IZLhs1xAm5SG5u84Rjzwd+89Hae3otgl5wvhLv
P43wfsacTadeJ4CmZY16qEHqqxC8P7sfay/b+w1YNNnLV6IMJTzTeNnne4+40Q96eafOHiI8Q9m7
3SSqOFoSq2mQlqKxn/YmHbju8/ObdGzulGjMjo/ywOeg3bQVx3w0egra168w9peDT6MnRDB4KTAc
KS+xsA3zje6BanKHqrTcaXO62vQUXAzzKKZ4rjoqcxxhHKY7b1reVEmSO5e7+UvVzXnRpnCeRL8u
IpsfDekJRaCSCv39QcZuBfQvjfxcI77tw7XzT+BxCmf8ZQW7fqkMzvMrNDqXRk6yqr8oOS0t+qyC
xH9tGAtvfcDlp6fYYR/jVY2dCffmwTemOsCLihfmC83fyWi7LNqPFW1YKU+kuLu9yQwLYlH68MWF
qXO13vsPMKSPVY8RwuH+VHAid3A0Ka2wrkhT0fJIjKRRdfM4SVZXyQ34pFziu5UbTHT73RNiedsL
cHqdKLGI5bHdVdKJkDW6FvvsFPJMEeAbLx/hBoMKl0oUZDB+gB9INmpyo6nd8BxuSV10qz0NLg71
kh4klaeLk1ykrPiyedJ5OWkoPmel/nSxkGp4fAGB+BTjAFq4s0qsVK6EFOvaY4k0lYy6veUfuIOA
brTHqqeOkT4OSYQeHz54+4AvieYYOLAsMl+43+J3hEsD3NSSkcrmRAS+sHZrNJ/jaGtyvlhiehgJ
s09ocEHYKh5iqOgIoUYRFJBClkvTq3b/wedVgHPwWbLudYhQVxGaEfVMsFh50qJbOmIZS+/t9CeN
CG72mSTknqELOEIkaIf32b8tatUcmJSA7A1DrlF9aKlOptVvcW1p6JPxpK5DHYKCHU438rquATg7
erKGRP2q/v7o18LDMLeUhGMRl6RM1ql6EqLEyouz0qD5yCyFBqMJ1JrxQ3m2n4OcZTpZzYC5jjYB
9Lo43qTYdTCbIZlNyvwL4/A8XlWN0mFOiAOETTvKc8XVd6vSgTVbKV3sTl9oGU3JAj6vsSBohCTS
VFpmiB6TnYN25yELHMtH8Sco4qJkn3Nkvsv0+U4t6iLp9W6P7LvAlsxJEr3g4ghygcpJj2aqDEbr
jTbfhLwsmLbUEZfI4lRbkJlounOefHi4XRFzBfQuy0ClfCBE4NJewQlLF0e23+KN0nf7rKZgH2K+
TjBH6PdMFz5M0mFFwbLSrWFchhv5PXJR0slBXkwfo93Y3Q095BvuXd3kQKdxmk8LxXYtjOliIyEF
Fk2uiUCXBk/3UpQQ70XuY0T6U+ir2PuRz2wB+IVXBhZ4TZ14WfHOB7hP6b7A0nQjb5w99agQnwRs
d4H1Eq9dR6a9GWsBvakWalOCqs9Qdv/b7ZnsWxMsRK36nwHQrcBF3AG7APTptEp1a0lm2tia2t3h
BvOc6B0TUcImLwfT91NY3OJVs3UV4weL1EWayhxawTCfT+SBlkyg97DW0kOEsqnknapgjg5T5YtN
gydnVwqq6RXen8lbOo49iVLIZm8SeBQPxuhh36BJH7cOTeoYpBn08xTFKKC5BiwuI62bQgR1SLXz
s8wMsuEEZjHEdTBk4FEkmZFqJ12RXKT7w9a7ENVx1i6c7Z6L8v2BWQW/LgKKDNS0VKuwynRmQvNv
PlH4vj9jIMu/z2g4yvIrVC2hsF07nldLyrAIH4PwWzPEOb63xTXlG/Yn3UWzl+XbeAyTHaRWz+CU
twg5EgbNOyO9ZGHkPPWIaerSKigplYmK7kszXQEEN9XOFky5EHIrqVdhl0cq9QYR+EwMqFHSczFP
kZjAZIo0BPOHIE1K3h6Gz9Bh8+9o121kOoPRPhPg52yutG+bOFu7mejzP5ewD5zKmMb/tA4+sxN6
BlQ1LZAhLbS3wx+MTIHLrPD/mG5QGsyFfukFDf8BFkGQIKgYgx5LdCBfpT82ke9c/i/vGo1ch+51
N+Yy78UWI4aOPAhw9+Yn/fe7JCXts2g3Sw+yzm3l+Fo/cLHYxBz3ijzWAsytH6vGSreZnsTrEE2s
LzNKvglKwtLVzjtdA67NU8OW8w68zNElLyIhLyQa/RZaedQB8uHkTBQf2PnAV228Ah0D+NJY3/y0
i53263AI+10Bj+CgsbUk7e+tBx0eTLekEPdF6lWMnuH/A/VyJiEA2MrX8Y1AUEeiHin/YV+wYuDT
gazTB72Osk0eQj6k08E1eHt4V0oY6ojEk6gVb8llCQhDJldNJQx+a4JTECZdD/zRNDLEEZZRzaXE
DGJBeEE3/GNWScg3ECCRoUKm/d4aTUZ76mpPIU32VKMlCtgzcNy95uK7+t45aotAza2mmRw8KzUv
UIJFZHsGzOf0K2Hkq/hlsf0WXBWIs8/S9SvC9eG5ThXrsTCdiR86YoAW6+Ttz0EZFyv007X/93y8
Ms7BwUpWV4Jul2hjDH4Vt9ibn/Y3KKjXe8qWR7vH4zKV/wUjOKZa2LjK8e83NxLY/Twdiih8cbFg
KKmOpUoaS+VOBxJQDX1QufO/z7Isb9roV5F5ZLJRsDW3/AddsorgmFCXvY9xZ2YaELUQTZUPSdgK
kQLSkZlUuRMgWVWGgXZSYtxjXsUu1ZEfJDwSfOlaJ1xMhUI0WIswner5PhBdFvY6DaTk36VgBb/W
lwOw+cygCaEO5D70TQoWyj+JPaMh6PK/y3sFicJRozRr3Q2rwNadcXMey3oDhM8L/FwkuLmxyrNP
mu8h7I8k1m6EciEP55BkLJhoOqmZj/1sJGfdgRCC7I96PpPr5bWydKTxaWGb1x4worVjGOPxS4mY
/eDA0HeQeswSE3dk/sQOofvWD6imLDZv3erb8Xx/SDg9KxTAn9FHIagyIcBsH/AERiPHsHyN1b2L
MQFgXyWFH6e0fhsDND97Qcuf1o4RojHME0MRSX+y1gCOznSo0lHUv8Q83pqk4gHK15kagjV03yxX
K6/Fson2AKL4fHbSiFcsqU+RBU6fQmv/2xPYA0OIQtJb3fXUDU5I17hOxVLDaR0MljB/LBT1BVCu
bR4n+vDKhKrbSdviHmCIiGVNzqbyLIIOstqhLnbQcdAKAqFH4imXUKHLyyE9KsibdfWq5X5SudxX
aDQgTUdtGdPI4SpAHCbMWclID8Zp3Pz+SiPywwPbTI9hGxzawednG58scLfvtDaWEcHfihR2f/J5
qhXmCDZzfsgmRGrW5oweRYz/HXlVRjgA17wApGdOje68tC4uAkaqfEDFr2IE+k+ZGbBo0MOcx54u
npAWq0BoQVKXtY7SDkN7tCIvMjaiJFQK18fo0aDSZtvqIPlrHvJUdvyC0/fN3oM2+GhY7bS99GGJ
6F33EmknY4nUB3BHnOvunshibr3o4ZNSfeSpqGpp1/i39xmxlUOFvNN1PKlIAAE5iQFVCNyFyei2
2DrT2A5lHcnw6GgRn2p2G2QCjzZoRYN9L/0UB6uwpYYnH9FUEo2UuLnCc82GMg47DzuJ0nZ4Jixe
qz1mJiCZN+CFUNUzSbG+aqjjA3hTf+H1aUeLjcS0slJ8Ln6iDmyT9JKV9UNV0hLQhmI0yJeE3+/8
KnvbBFOqjBqhyZ7x9PVCfy419e2ZWtf30hgl9VWs5lRzR65I9Ardtw4B2GAzTlapMNfdpZGHGUaj
2CoztxwD61n0+a94a+2q9wK/5b8kCqJ8vtqYJ7SHGB4FeuRkMIfblyZrSko0gbD209q6eVKjJTz1
glfnERa5Fw5NiOqQivplvhUVZY4EaipXK9GQoEnbcEIJVEZ+YYKt23vdILKu+FrOSQjK6CSsfIll
mvyCFBQ1OGzxvfcS2dvdVghekiT/MGLhOCin/M0fAOE5OBcV5LFSGRfqtj3b4R36WJKB6dc/bcLN
k+7m1xy0PmxddjuDL0F0/wBPwH67Pl3w8T0WEMPGoV+BPL4v1hmGhOwgixIB/wR5NfC1iyZQ+3/1
iAoswvQDa9TkCS/q99njZG+8dGMlMEWDzgmV2FiinD5iy83g3VX4fxNH5lP16l3PFMBuKzhVP5JO
eLgp3CZsfIWmm9SD6ag0bGMUD182tP1G2KuSXTyuLOciSBGsqscmyrGkiXFqJtrEHvCyOn463vjO
0Rnv8mdLISSE0cyisnDAxjkYnWqeBtILPtpZjH7p+J/PGrm2CLa5ofZSfa+AO5zFohp+G8aTpnDm
GAK7CU1Lj8UQEc5G8RRn0SuelF32Gwf0ehn7uKFzhEADqbvOXYWIQsnvTtnvMazbdtrbhDl0lvU6
OMH58n7+Z/GlK7Q0CJzsUPjf04HHe7T5uh+7rjYJa5ngTajqmrM+gmhUXjgXRWmPyM+ZUzzJHI+U
2GZFnxNwCJu/SCh7wkrUK1ZaKn4zwnw7Gx+BwboRXoCBX6vJVM9i5lIUgxe7FXIOVe/XThc/PSmg
pM/iXXqufL95mIIMHdEH1r3KUpOVbX/lqMzvc758159/sOwjf2B5vr/u3NOQsgiYcpCi4pyw4iTU
ZOaUHnpUBoJoDUURTfT4/lnsW5kaLc2Txs0grCLu8aLFbzuGISMxBOs+WatJi9LjRVeNZIFlDMzC
F2/dPa8q9vO3BuL9A8nCd15ZHuQTSzjKbNoVVPDIMOXkshGoxDas2nEQcLc7Qlec3vCstIe6xtOt
RaxMlKzLSrUJEeCbsrzcyRg/GeJiAXcGq2GE5dtaGSft06mt2KChEjrHLy0IfU7w3pyHw5lTktSX
EoDTkWirPHxvME0O+wzNo0o7U1Hu5kjSzWHGuHlZH3IAU19Hd05qVmmL6Z7I9Xb7O3ew+mRF/IUe
Y/pvTBp8cbh5Wszofz+R1sldg0Trm61zxPDGPYjePqObzh67Z+UCZOCuGLJEUHNxoRr6CvdACiJc
RTWVpNBGfWI6zfuqkPco39voHuA3hZxH5ELP/y5EMPt95gms7IDsZ+7mGL9BouIx0p3pGi7HR1Bt
UJs2vc+VH1wBu2vYovUkpVR8oK48V24mfaSThhEHr1y5l7ksrMYi7pea7pMsDN8RCGIR0iFv39Zl
tCMgOZAabr47ZdFtiJdH2w6OHdxXfvvEL+a6Mm2bLNy2r/tfIntwp3DW6P5aqPJhIx/4fzMe1P+B
bJRw99/OdZrz+tiC2x5/kfsp2I8Og6kM7N7TLqnQvkB/2nkvJDYvpa+5cv7DOjpLMBpx17Betmwm
PU1Q0IBuMDWa4aUcHe8GIARga4I4QjyQs+iHOOeI+WxO2jrQKb2Xw/DuXt+3AMZ/i9a239YHabMH
9tsy3ahKYCLqJ8EB/6rv3Z5xN2tCQe17lJsr6I/oNRqCNnWAxGVPYKD2n8bdrR0gzQZ7k9lG9/Fd
/31IYa2E0pvkO+f6422Hr11WJ8twjNwgLdDLUbGT/yQOLjN92f2yfivPilUBdsh71DxYASBsloW7
aghiHnnEbvwXTsTuonxdO7yHvMfFdI5CxIac3Qs2CtmduRxZQRXfp6ZZVix/mver1udtOwZEFwwq
/06Pep5wMhIvAObXpD4rzrq5h2Qi0+hxMRhe0EnE3MzSWED/DtEvMjHXC3q6RruWLCYAMKagRZC0
Uw03quQtSlENLJJlMIKPeyh6NcS51JLLwIh3Jc/B4xDMoNzetJfVOZM/1BgIbl+2ywtORZ3zgHrY
LbIaJ4oQmcofIZ3ueSN5231z+PnT5xk779JhUqgmziGjfpbCtQvCmYHWZ5kZzEE1IdzaQg4idnJZ
JOslGbnKHRjerk84zaZwVFic9sBKg7N0cQhRYhkBQ8ZcI3nFn4sWR0JkhAsSRM6L24uxtBu00e/k
WBwjFB7GY28nzhCFvp98nfDB4O/c06ueVKJSBsAh+WHebEmJsm56NEab+uQAfBXDkho41YkDXFcT
Ih9sELsvsZPN1OrDGtQ4NcUTDAnHuaBHWeHYaCNvJpy6E1PvCwOfXoipv81KQpVEMyX2hjG/OyMT
1XiKYx8/N/spQrj0+XWI5/7GyST7NLaMhxur0Fu6AwLTp9RC7nsTfc3OG81JhVn9epLIz8E11hca
ByOIjj4yhTup4XgFdC49fGngBZZEcdPqXjRUG6ezTcS4ntdjtFG0H8yh5zsJEh8pXDk1R+zBcSaV
IThMTx+X7jbZMd9n8Ii/C8fS+vBp6mybLBgcOnkcyqReLAgvIgPsWiLr0kedVq0RQ3zUk9GlHJg5
WLEyDO7VJ59fhG2Y7aAHu5qDvOABcwOBkmnXCatx8r5+h1CD8iSIoalfzV9i8bSBjMTJHLBDBVQW
gvdZKJW/oNRESkXQnxgTlU8etxe45443Nig5QnuhBQqm2QiVb2Ut5eCQzPdUI8sHB6QGm1WD3doj
tys/nqqvgAytRs1bX+DkesvEl76LPZXLfso3CEUrkd+IoxfsOJtNv/6m4nOk/hKEONHe03FhYfPg
3m6BgUIpVbJUcI49UKaM18uITkVy7KEsU7GBYRN69PYXpJrqhWdAIX55TUwb5ls/fRy8/Pu0t+Qj
1+Es36efpQWvTzj2mHjzluYNTdxDES8YMbfWPaCxA7Po5dxXgJrI8xfoIhUDMrTifWcY3jZG0IYH
jcBe9ju8fykXGfxaa6/G9ycgA99ZqlysrrcuKnJrO748LWl6mDnxfHtiuZbEX7AagV4xb9z0Kjtw
uX1cU5oDPLDtPQvXP9i4RfeqyIGjAfvhWWymnHl/0MMvwpR+uqsGfLVfwh+Y0EfAIBgck3oJnt92
ZYaihDvEFBpqDZJ4y7+4SsGop2QGsL/pwJITz3ka5b5J6WF1wKv9o01lYYyIav8Qecx8jqKOja09
pvy7xUeNOMrtBT3351nCkNIQO/I08QBewGGzy//bUEdMkGw7Z0sdNEcGJPH8PCk/MTZkV9vD4OgL
duMLwJcEt3ISsYZa8dfwLmvOLSw5GLGkGeN3qNdskbJDVQ7cFbK4jLM2cluAa2B3eHzU7evNJI7t
aHATZryi7ZtCGQPN5TtBL07gHCwW0+mS+KPHGXaT+e1Sh5sbayLmqVG/UBtxEJvZrMA2aFLztYsj
Z2cn4yMFhYca59P9uvul7VDnnPjDxacACR7DTQECugLRS9PN1CEVTyegUO2gmTB6SGJ50v0UhMv1
fnNQp+bjcVDufAUSrrCrgK+YYbF/prJpI0dceQs9QbDwGbsohNu6abrpN3tXnzyQ/dTe49zKzowt
qoAd874/ODdjebooVHNaxemeQ3hxspalYbso4PHaj6U2Fvj9co2sGBLzXJObmBlImpa05S1lukLk
eadPT/C+LnnE7RZ9GnmfmifGrEcvPVp4dJ5AL1h9drhJmwjiV6tV6YeKEVtnpnBSC5G3KFZnLyCF
geZv2Tzur+XffheQXlnLUrv9q8IPjOOnyN2uW08gmD93BU8l8bX+mhm5TK76Y3dgFOaxk/aXVdJ5
FtJQpTmquUg/3MGfgDL9vb8d14rC7Q8Uw+1SNQ+QXsrwRZnuVw16wowpUJXkDJsWI8wePhqX4ZHv
huLrERz9X9aMygNNKqcwAaJar576OqM7nHLWKnVOpJhNDHCVFfqS3Ml7scYYq42mJqUfLS9BEJu6
beGnSqUPjgNke5V2RuXPtaqQ1574PtnlcjjPl8AzDoLLGNT5cvZkbLFYpkVlvZtIKjH81uY0W15Q
SB7hUN2PODXVtY228PxgX40saqRyksZ5uJ7tcbA0enOv6dvrlrttknmTXGc1NTdcFsc+DyYKyldL
um66cYqWHrssOuMfyBi2d1fkT25TfvyQRTK4yVZfPq60o7Swgbeccd5CtMJJ1N+vsOH5U88OEwoM
JtSYx7yCvAUpbnJqh4QUMp6HeZSJ8K24hRyPA8dO6Epr3juuu3psb3UoRkVU/7TZ7ink8qwEhnnX
W3J8HyJ1Sa0vk7cC4sbuERUi+SXI/aamBNH70ulrdkq4FBIpG+yhlYJCs+1O/s4GWTg7kxDjEGiK
P0g3FqEt78h3H2RMTM0/b2domiF/5Bp6kyAqdEpoBsvwtnN2/L6No9xVMi0+naQQ+Bpve8hhsNKi
yxQTs9zB86W6Onyxe1bDEJy6qBB4fXa19XfV7vQwR03TixxGSdgh0Tdah/YFNcKg0KyQfz/EMHIM
yRtJfWIfAp6YlDyw2PO07NuWSxJrWXrF9n4qtLxwNRpR3AbNpzJ6TRRYKoB/BS8HvroTVUeHEVVV
cqzDqV+M3nQvbtULLVdflKQrzRhABctaxaCL7G3WOWDsKV0t1Hx2Hnu8xnopLdkZ+sQLJZwl8Ptk
o3kLoHzGDRQcJklgGi8cf/Il1ul8KjofCN9ogcg6Qb6QxweOdrZXD/vsF5EECUa9Xm51uKiR9OaW
3bqhE4iLZ7c+uqCr/fk8EVnuOmIg5yNcFlel341Xx6pKlRwvrZZIoHy9BiNnpx7REHvRXA+GsX/J
xAp5J5EA7avDPsBxMYnxqq96b6rYJJEU4Dv8x1tL0G5rGFqSoZ+/3nSja31rnQ/xKli+zGEmhKae
fgyPQpPiNsVZkXqRYS1b9HbjIe27bJhw4Xb3bMhblKENIgPuwdJvU7YOh2UoXdDyTtoZqBJRiGDG
kqPQhEeI5zs7umywbnBE3s3u/TV3H27Ttb8WnYiQlTfUklRpRuNovf5+JnHKkZcQhA3kWQh1LIck
mCfb7Wusse4zxFzixu+peca66cKAg+npOvLsHrUo0uxdbN4MrwXZ9nwj7RYWj4+OYc77rBmJfV3i
3QRcZEZaJmr6Qz5f2wObMX4C2dFqhorQMiKAjmAxh1XotAoYyxHlMuy1vIu/nCRzJJ56x5g4vn9a
iydNDC/vmedd7xtPGM0rGEczmmwDrzru7lwyl4oARysA1ms4qwfw/wXTOYvneXsekJTz6py/WUL9
QlWbO3rLcWeGRW3Nna2mSck530fRpV4D4AWWzQdlozbJgiJr2yKcWaBsSp3kw2f8wmZ6IkjIYpLF
rdx7xkmoBG8ClUtVbW5/Bj1XmqZJ3rgw6b1fwntA8a5uhsPEH1UvfZkMOHKa50aR1mv19sUumT76
DaxZYsMqbuCLqXkofAA+ugj1zMQabh1DgfjebI88kLNNF0FXn/lTYWXHdb/nU6NspXgCUHci0Y+G
vAC6Jz1jVweIUau9sw7q1qr+pKRB/Nb9PUKYJtowVwwBmdxpbAZMkfsOl6RtcF1cba46IQuvdKZU
FPNOE5D494D1vuCG3K4DvMd4dTFBAuRvV93te6zTd+G18oRFPMylM2AcFkInKalQJ1zBNoxavYnl
UJ288UzOrjsN4NMQFjw2bjubxE4Q4ud16cDtUeGOExm2kTSdj+jcSjLsbMK06yTyMZhgpSflZTWA
ZUl+LR5MOYdb7dX658TUuHET83u4QjTDG0vBFqTBGMFecAh2VR5IvbXarPPPKDUMlyTmtUScJqzt
CmHuM1esRdJaztCtbghOvg0ByVYYDRIx2RzZRraputFpqQAGlQiOSBaidRIRsTO/S0tN1AkjClYn
3uBEAonxUkX6Thz9ebfmnHKZG7CohhYQJurQ36hJZ31sAhkJje12bVeBNIK418NjnvZCMnuhlADM
Jq9AFQaWjs0pv193WR33stIgVFfUW7MPwiK3dN9UmGK4g6ZmAHD3zP9nOfezCExO+YXfVn3bkvXB
AKFbGZOtJzfyAlzbcL//ToQUDRVUawV0fkRoWlN0HJ1NaJ3lT2zJ6lEmdRy82JdxI57D9sNjzRQp
vhW1+CIHLCAPIlQ4uiDyvRBN0lIt5EidxTL30/fSO0dSGrVLHIf5lsJQI20Ze+l1LNHml4/f1Z+B
3UNKOZ6JpnuScgHS1mOgKHhNCdVIxk3h9ZTw13o4iWOKZdCcqTTPkB7/KSfL6Sc9EMXYkkUQ1oQ+
JWuIbI3UClarUPkGMKT0frGlymdjKqLrh/eoNA0OgsAHqwjrXU4DBpjuvpLuK/9OY2v4I0uNhyKN
2oMER4N0bHFMvo/MlaUtpZUlUixPH76O3mwV2Oh5b4KpfLoBVPzkZ+PEHb6K3+Fv4p7l5ucbeJFL
ANsYoFQmplez546gX8nPXifGr52d8Xt1McTkYtuErLwtb+/zt0Mynu81bPJejn77sFvEMHAbDRFl
NSMyR3hbox2mBja4gQ6Q5tlf+USIayFPNV/g0L6Dzg3dmKvzSCDZamv96HRRFzsu36TDjOoRiMc7
rDE9SuaTRGFW7B4S7Ilnjkg8eeNuKKLSJETwo+5932FDgB1WzGmDeosg/TpNQHQJ12fmD061GSF1
HEn8/zNIE9Rp/dQLxPYner0v+ndHsWYRSOjnmDay7YDbX86XieZO57xigjUnR1bed/8qMRMAJwon
Z7tdPj0ySApNiCzXP7mybbAG475Z8Ax5iO/s85JRYiyArAvkLLWeYTLS+VbJIPXjj+pykW2Afi5P
PflQgWyVhoglVRtyqeOYbdVWBQ5K8K+iyqCn7Cc5FnonC5cTplppbsdtZmCmTsMzInk2RQE1zCfq
8sULtEDHcn3R1Rbkr7CKMAMf44A6JnLs342eq3798rsdRiT6j84hoBWACQpcyXSQBK3axu5+Nzop
W0cV9ttk7cITuRg/Fk6kwaU+zDF8pgoQBVeNY+l/qKO1QuO3VgQiCuKCHYslTapwUhjPbpPjjc2t
DaTOPwphzP6h78qeg00BfW6R3ZE5F3EUIKBY/F3WX7sWWzrUrbf05csVaYJxQRxxkAZe9H3hVIlE
XOe+C1aPr+8Ib4/TeVSGbK3mGwM2mpH+D4IvKUGXfOkTUa5UYjGGkQnRo6kz78zAaq1/MKMnJGDR
IS3etQEKGdYeBpHPlqXUUTokcJjyxZyH2zCQ9X+6Vrs7fO2JFbNJ8UeQuDru+Td3CP2PLw+YZjrV
6MQbSq0nt+W4u1XY/mBgkq06fpcZLokZRvtti8/fyNIvGqUZ0u01f2szX40biQdl+BIeFgOQbc7M
yD6Y/xw9mP6AOU2H2qfKd195wuP3LGdU8X00y6upLESo2k2Eonm0v3mHRdSbmkpIFjPDVKV5RLOY
G20EfyPm0hUjLRtnfk8fhvRzzVHuEavTGCuV1GZfGypToRHgw3WSYzbSOZ+6Mrr8T+GwpccpIWZ0
YilUrfdyVphBN8uXUZLLEVKsboqfrHiPJ+kf0ZdrIv/lgpJNHuNuX+yeDmN2EW+wM2VFPppkD+LI
LdJpVzCRThzcrZzLccHnvcksHhXsWgMzBWb8V0n5ukg4HABPaD/GJad580AQGs4MRePSIxK3uccs
rFXiS2wkMDq3PzMhf12OhHu2xnC/xBvMUaQjLv76yEOp629YmIl2s7C3DJqRjM0aC1ESNzpdaRPA
uc8QUfh9QKyG2i0iwl1hBt7oIvdYgif06PP65BisOHk7pGQ1Fbb+Zhjk7Rbk2zMzK0JjHPZv2R+Y
+wIeJwYCa69HdJEgKUezYueTfJ6rz8F+GsQCX2jfCkZC5bLF1TsjSiFk9EpahYnKFpq7h4HJhj51
Taqwx515QvJSzrb8ch8hZQc829h4EVwGRota7fasrb4vp4VDDOJDq9Pmhkmu90Yol2hBDTgWQZVb
vEUkXSBvVcaUOc6EKOC3nhvOrXJWhYafHbUNi0aQmDwdEsI9W8fx/XaRjEpuN8GQQUdzLYW4F9YW
FcKJZH+5UUI+gxpHv1oPyB01xUWO9mT9KFoC44Dln1KXOD8+UKOUfU0v9HGdpCYIcmh/uSebYlw2
4Iy7KjIwWOwUWjoGcT7vK8kEQU1qwJn0EzvsPHGzHshrzZZW5JWNA9CRA8Aumdz8ewTWAzqqkSZh
Mv4loJ5jGxUBaOjpljkoX8sGEnOwQL2ToKpW6hSa0om79l71VJz3eh8/M4J1vK7Lm+N7b5Oxsrov
PiezNjwdfkVeQgXY+7qlanH73+EBynU78r5fHs6QFUUg8AJKMN5Jy1dDrtJWPgI/7Lvqn8j5cOpE
zEcd+ePpSfHWgj/84n0qxOy33RBduFqI4mRPInIhx9188tNb2CR8mY+13PVMRYaiZV0kb92jW4P/
dSz1yXp290xMjjMcJ9CYMTykeqXSjRX7hVDHsAGAHrO0Y0qP625gsB45ismEaw3qs92u1eVYCrvY
jJ1r+npXnaaVUHFZDM5ZBF3BwFViOerR8YEd4Z0kaHM4vATgIMmZDA2sVn6/xyWkTTt6KNihKiGx
aGQFv6QwkRd3oDjgTklO/lOW/Rryi3LUxz2/KjD604bckGaYHTTflgcKw8Qqqrj06lw8YKnU7AYc
029nG/F42oMwnXzEDIQMVEy1MbZJNTxyn53vHSg8PrjufQbw1FTu2thTzeXpCgx0LAVyzY37153Q
fY5epoWOxAiX/37P9WuG48fr3bsRK97ldNCq1mELLJsLeYxYH6H1ai5VjiYggyjno9EyZRvNSmNh
z/PhjzhkFY/NVg+ygmlLA8yOvHJS+z+UADu+gp7FIUzmvlzhNoVJvACRndd1QtQXKudRUDXPE04H
aNtsUEvFt+tP72OFFwynz8RbP8vpC4fKNTsEg0L8MK2a1gDd+OW4Jw7oJ3i/pt1vtWisWKiIk4pi
5Dhny+2Re9gBBe6YWegrnVZFPgjnUk8iz8Pm0ufaq0o9bg+t293PgzdAKt3Vx4u8Z/N2VtCUnHQF
k/LmduThMODwZULRWLIlthEpeyNaKUQ4JA7tiXn7jMeurQIES+oOyyPts0iXyJ7C+OFY8Nq+k6/B
koWY61TCw0U1Jz8ESMzouPUSArr/gV30VuYzGbSzvqoBKgex24KIjBQm1MluyVHPcwGX9RpF1FEO
GR9nWXCtaCDh3hJu2PHxiLj4YdGFDNo4sEgae8uBlGLc7gxsEZU5662bLsltnSWvzRDIUNtCLvLF
/maA7rtYNMwUGoIipL3WCgDEt3MKXkkNRZZooqSnTCZBQjjKwbF9RSiDdXEN3f92sBEnlUFMMr/r
rvKpBi2P1OqSWauTZrHVrS+Me6ZvkOh2e8AF6aP/aTMruWkC6awSKZwclQZwR6GjJVJhjyAK/d59
Qn5pIIo6vuGAMkJX2vEFwX77N9vScZPIl8TwpXmsYRpkbal8FYMiRP3NCyR350zIAaE78NVauL9U
ZEJOjcKwbrmuTGUYOcI0esZPpcFdcalBZxcZB4fpCAijICF3dEkatfNPTejG9p/UKkMxFUa0QWy6
FUMPfYrqsXwxZooVN2vrQcJ43pKpFe4YhIoCztGOCoY7Dhnt6ccpPqv+3NgHwu3s3sGhH5cofA4M
P0y1jP/oUVlpjEbpqZ+BgkfbbamNy/fl/j8yMChPnsgddwMbYNYJeNBhoRhz9TNr9ChC2PvnAZXG
j2/q56B75M0cGnK+FvxoZiKo3Zp5JNjp2bFKwFH0Zsgqc2i8L92XLBETEsX2eZ/hbgtIUXZONlSF
p6xUmZ4/BCZr2+dB/iXz42AD3RF5LIcU+9rKmFhrfsSfJLGEQhOPQm/q7YDVvQjgDQbymG1Hd07a
agwBbFT2X2UqaEWhNpXnnhKwUaLjgHaCb1KrHSgUQD5Jc39rco8utVoLJ5XB8Wdy245D6PbrG2ws
dLXr3rWpSv04UAaKUTDVF/QcwDpoRVnIUBgTZ3+oExZnSgmp1pobbRIsOgX4XLRPVrk7X8xGlsin
X65R1/6aZtEjk+edi9vutt5Jwo55V72tvxUdwgcuHflqAS8islop8OLRteAZlpXmgF0hDga3C5YO
7mmD1qhRT9556uRW4IFhrLZquufkTPRYX8nyzgSgImN1g+zeabsGXLl6Is6UrAGT2WZp2uJS7Eyx
RYUiwhBLweTfGdxryYvveEP7OXt8tJF720iNP7YEddne7io0G4TbPmiPOUdK78ievdM9r4kEM9C6
LoPs7JCgQXVhVG2NnfBJ+1aDqhkiZoeE+4lo6iivZPmq+xJinBQ/0l+z7K5/y9oa6MyrfYZpyiUQ
cZWG+/9hkfqWlRCwIRaelm6Rt1BUlCx8tj4RXj6lHoHzt5Ly+92LCh/PvnzwkLgPPuSpmaVFT8kp
ojbEwP6nJBjJ/IRZVxfE+sDmYuIPwfmoXXfEOiOx/DleTmYUJLPW2009GpcKiuZPKX4yv+UoUuFE
1HVXMUDFsTwxPiR4yuQvdatxwE7QbG1294IjDm/pv4Kj4di3JdNochIG/XZUEbgb3xZ+Adhu17pH
p1d997Shjzhi8UiFJNn2RZ8xzgTgo/z8HXRDjA3d1KRiYqTf8rnPy09h7V4ONW2itDol0eRLAJ6d
fwsFwZ66OxaUiCI/tm05046e+1ToG1Y5EGqiT6pR6HxYmmo9GsLS28128sdRb1DVm2ZOlQjEICby
QR1a9OJiH2GG17lzCQTW4J5N4Wbzt1xj92VJ866mLsMHypVUwD3xsvEz4ZV16N4qjFxOPsKHtR4s
2vavHksSJAxXvPqK1Ldcf8d5She64Z8XVcBdH675pWTFPyyKMEO6kXkZf0J+3ZwmM7qk1jjVYnMk
HCOhONvYCm4jlE95+tL1Mjue9QewCJyEqcHjvieYMZKAK2IAW6tNa5iia2n5Pc7jtJj0HhUVfl9H
u8cDOlhtWsKNWcXbNA8ujgnHYOnuOmv/3aE8i5qWHt98/3sBRZ9u9apRd9LzsVNN4S4EyHrq0UHi
Gj1aDHqU3bHyy3cwNAMXoz2bDLVYgxN4H9d0sU6zWgiNDmncmhPhUos9ybOcUnkjFAK+LT8zrPH6
eDEkNsQ3J6FvS1DWOoMeSGAdnBAH8s6a3rxJVxV2eewM7twXamWHYmkpIyccqTu6LyGlfY82d3cD
VP3O9iV6DqkpUG3+GPqJvmS0D0xpiSZB6A/ljpzgZVXqBmrxIus7U3U1mz6M9im2+LxLn5pzklNy
Z5XtL6LjRJz6TCEMUkm2aWJcRm5ontvaVrEiqQ/ilvPEuVMXWgJ0Eo1nr0FUBAJaeEo3Oprq7VIb
jUbffQ59L/7ne+axeBis/TdJxpbeC5hcIyPpDPbwUt2rROIZr6Ikb8TuIY8pC6RrdMVsHe7K8V06
JCaNP8gNPseUNrJXe8N5xIoAfAmFRuDUfqLZ1zb/AE+/6dIjidKfrXrwvRCELC3Eohf073ySdNYv
dMsxeHtMv6REjitKUk750CWB6vfMZHcDgJcTV9Fe9SvvnropAW3Ely0E4lBF6nbUcQx1ley14fH0
/FdKY7vfZ+rj6ngbIUp+JuQdhM4Txzbw6gsIITWJCYN8ymd0/gEZXoYd5DsKXzl1KaN39z7C7L7v
srWc5I3t7m7opYNTkttU62zUEZdSnpK9SJr1MI0ZU8vbw9he4i8Kw+lW++Mg3Yee7SfW4y9okFWz
IQoGsDVm10KZ/0CyQ0uDPI4d4KFYcWjZkHRyKX4mh6v4jfmIaCA8TyJBDvRjMxbJo+nNRuH7ca5p
fnckJZVM4GoiRJwtlyVaEZw0cS4dUZsKFJx09FVCwTqncxQVfNCOEkzfpucHUf/noRRSngFAi9gu
MkDvOMHkG2mESVL35X632iE0LQCcBMXAyyluhSO4dGLdu+EvCysksY2yuoZjk6pPWRbEemeQQBTV
tIayt/IgWS4JnwPPf5nDA1SN9n2bKJGA3yKvXyxkv1pulI/sLoKLkXiuc9Ff+lJe+EZKoAb1mEYa
oXz4yXqncElDk+rA/9vnx2ZUCRfdg3uMSyhsFs8c7aQ5NvuU7Gyrp8j/TCtc1jAed8K6m+pAgzUK
bojCUrWL5XxqZHjEunPDywUHnxEm7X4Vb/CXl9nw2xvSdONi4xEHPB/9jXHfcfR4kViP3r9veScz
9ra18XYjy+dZV+8PxYRfYzK5cHfK3INFX78P67ciOdpIaa/EH9+7q6xe5fJmjhFXZgAmVWPiZwJe
8WKHWzHrrVsYu8r7dwIGXcttFZRNGrAeHtQoZe8IjTutOPTCrF6ozEUL/59Rz7VOj1Jg98qFluMK
HSWOCvCGySJmA/6p0JyuH6Gn4QSCiRM9FkfOnv3DkTGyGSIe8SP0s0xOOoXrw4lOEg454cy+yZu7
WJwtzKVUBQCbhKwo0q6A70e/pJSmrcKGbUH7DnRGYXW7YpCoHu+j9Mh74kJ5y5pBqfpfsDret2qf
IGJnTH1qzkRDpR4EPJ6UbRgrVLH/K4cDLZMx9z+tJg5qvOD2S6TWcTvTrZ7aOadn/UeiYja2f8HE
XNXQhvcHHmKN/Cc1jbU01IZis/fbYwXVQy7lKnVT1zgTellXEa1jR5XJbeXXnoJst7EpCPDpA2kI
k7aoHiJWEH86JFBV5m8hDvRPLtNZNfJzvh254dnXo0pP4xU6ZTYU+eOiloHsJaoYlwee0HOuIJeQ
EmyeCtSqmU3k0F8ruc7+C+F0HKO3CIwTuJyMjyUGzwZET8EAQ9TXZIQcTIWkSqcMkMue6h7iR9g/
yc+4hgn4F7kTRCMHWRTZf+tI0UznUgQDr64QQjGJJ1zqHY8LAVWEry57ZKFkrqn1aY9YuOuRiaWh
tIIq5HUy0d1uLOxPG4FpHLjIGi4op5S1lRHOYXUmjy7pJlRn0U9M+hUi7EPfsCR84+aM0hx6dMQw
+00ptjxxZ5P9QlVSaUjZHMpTO7QctayHPy6BnjqzCsm5PNY3xFrGSu+G35kLHMHceLylrNgGpgpf
7MQaXGpg0v50VexzLB4hwL9BMJ0gNd8P634t4xTz/MEWl8Mtu3BrM1A3CWYVC3pe8VwcvOa2+pdY
LBL52hwjwtZz/0YM9CqDH556UBXuCNY+iy8nzZBZR8moDQQEMcPDjFvrORyD0LJy1Wtvl9abhcxf
zN1Ni7mMnh79SbMNa4T9n9GUIJSmFZ0bTJvDxPQ6M/5O7e5CUxVtVMioF+9FBvHOq7NBC2nyvsy6
0AzETLAQsTjBi7lMTWsXzlPa72L7WMFxkRbwvSOrcK11+FlpAW6P+jSDQYH8MpeQ1bIEJqoqBTen
7BsWIYP/lmWgcXEur7oIu7vzF7IslWWhv91+SUtUBeFWeBvPI0dTpKSPEXBttqDK6a2GyDd4XVBa
HCL3GRBL7QH8nWH/ld+egDdJfx0x5s+/OLD7TgLmrYlK6mTu/8KrcBJTlzd6N6j/41aPOXMAT401
uZsrdbJulLohnQEJaOgeMEPhB6k6uxxY88zn53gz9zqMMpn0xJYlbJCrODX5QciH1wurSB9mFB27
1rY+CPPANQLpy1j7D3+V7aJ7dnqH6gIOMW45edv7bfC7s5y0gfc/oHogSBhiirNdSm6f4S61w/1k
4qJivIjvcP92nb/Ag/duKo8JdO9T0AfZnlBph0LnIf71wCsv9MOsy5+jDdU0KyaK3XuvDYwhtw8y
QsIwmDXMwUDutJ/5xYyV0OX6D+avU1HWuf+0bP2e6kbWFkgC3b7cUbApGrTLfFTlKunZGnUo4cmu
mskI+cFWPYf8Xzk1jWJoMwJ3FGr72E+y1dhiVQeRNgYlqzqx4LnBPk0iIGAxMMvTeLBNcPt9NTSS
eKAZ17A/9pen8+QtXTESMFIvkDG4CDQqMn5w0HY2OMFli4JiIfwbww276TPK5Gc2kYjFMRfFsQD+
xxWQR7m04YLI3ojDwG2oxE0eytNjm/g3ll2Rd2bYhKYA3RNs6L6nbSMwteBZuWkjVvNdgTxaD8uY
ApAeFjYSDV5zj7TU/lTa/1myGuEsTpYMX0CaOrSfyHcLUUnIFchnzjonVW++18Gp4r2EbDoJFF+R
/HGvtR3ckG0KvI6A03O5F5FbPBFaRdXg1uolkwBcl4XU7i06UVLJtoj4/aGLv94luvAMXMF3SAXt
EpDzlS/QX5qRjMaNlFwChdj/Z1lSd9JaHtP8oWJ97MLd0FTV+7IX+GEFDqvkrEoAVPAnLECiFW5X
Jy733quUco3F0QvOeXmMOKwOw92iBX6+z8BrZJYOEE3r5P3LeAh8lfweDqF+5o42iQwtZBBrGzf8
HDqAWXDl/Uyg25/1HcyD1YrhNutjwlPRSgp2mFHn7BaNZ7hgQt3t/ZTheQ69k3SwcQBWmPs8RTPn
5zNw5msQ1bvp2Nt+2lczF/40Qk5dHGxGBEL/moQJH91WVtbhAf3EbJDyOYiJjAajixpuOpysgn3S
zg05mlErCl+qJkQJfnsh4qcckoRmeUVeqHwue8z7Ezq5U/PEby0G57KoOYjLNcM0VZUFEqTzQexv
k55u/N+yTLntH9UcPCek6AnuB5JHmAs0tqFasS5O/MZ3LcEWejU2kAZKgYS6C0AXMnK8DaecNj0J
6NtTNquFo+s+yzwVVGgRe5UT7RsGE8PM9UKlCAszD1bL4jVsbhcAo8qjAzuVJ8pmcfDCk9Uy75Zx
Rae6tW6wDY9DSVpaXPJw7kdosdTUoayqNGphLq+3LKvJTply7mauQ69g2aXDOwELvGmaPJzYPsry
NqiJQlK4nZgqtiX8gHDy+gBlcTHis9hMQ2KgIcZx7hFgzzGa0SUHZ4W4iSDzti5nf3sK+GBL2OHe
tOlN3gw0F65pAHFwt1TTPIgSzgxEArJgvInlNamPB3RUsw5K1PsNv8DMs9DmmyAPmHAUFk7WjRFr
cX1ZK++H032/XzLGbns1bsXSbhy+sAFVOM8dGvC8SpYMQLl2SN8lVHCExKVUiLRMnf1vkq0r4Zrs
WNHqwkrtasl8hiU3j7Z+9V6NV/4TJWXMM9R2X6sXqJZsVHpm/fy9O5fzRLZyEb6pT6PEprtGlJUN
DycBe2UrElZKkzRjJ2rIA3jLvLRvaY67sJU2+t4wUU+wlfOAw0rRV0sBv4iFJiy8j3zE3Q43f6XP
kRYqOPvnvKDMWuwWFxTF9A164b5S35tb9pE5MG6OhJUIt8VzsPfgcCAtVva/TPDLxT1HWx17QFP9
hzexHJO1ZA+mV2oEPOsizixfkQYL+YVGZb+abEpIZaBHGGR/b4cGFAHEgJbO6AzNg7WlAqoUTbl0
aU01b9i0VINayxq+O6QvZH01LNXAdWMVKpErnjrbl+yJU5AM3dVQ2hFKmlXSqWEarf4sV51AwoP9
N0pR94jxkxmCpmAW4An7TDYH/NREAZIjy23QPZVjXnnLQglSiTG9G3BXT7thZGeE5zPVyQxZsO4R
elNonoAmSnDyC6gQslYrV4Cl3Sm2blSvY3mN9dnIta+6YxvJKa709O/+uh+qO0aXRR3vawP4Z1Lg
h/wGHLzlChezcXovogm6+GJ+2+vY9cf8OtYsaYAT8N2oKIXwcGV28YEPcIsQQyj0pCtSd7mGLYcD
I/pn3InpdXYJTmkMEJtlRBNOrs4NqqBGnJXUT8eWCvNqK3zwcI7oi7lrePDJrjE+EXrfN6Pb9Uzg
ew8aIRmfgarMb4CRyaKZtl0JDRZ0uZvpRKbS7pZe3IIMyO1Zp54MphVP485H1812nTG664hDK55o
BlG3ya5tLvvo63jZVMkwPgWbDRrB4DQuvD3Rx33/ciaCouklAkQROer63SV0xnfoshsbbWwC/L51
T883AEDMgycskusjwApunRweJ7VkxcnLajqa963bX1jarjDGBaH4WYGp40AiBgdDo9+ezfnXpJOw
06veK3Ki2t37TedIRk+6Xc45HQbCgo07cUey91K8evq/Z1JrJVYUxTcXhBj7zBBJSIsBkxrjgf+G
wIuBqOsraZo+N4kqvR/dVHabTRWP/4hMmJ8M4tDXe/59tvhIRks2D+GYB6LYSXg3tickf2yELgQX
dkW+7Gm38PamX7LECNQo6gTwJ83wBQAyNOo9AN1nOGmiJxzEPnDjJauPv3CQ6yv1uM/0tet5S4FT
ywpMqNj4OvfACZrUXXSY0PPYG7aE18B20L+BRA507qHfRWg1Joseg2ASZrKVXXeXEAiekrOBaveU
hB64CT4C73xNIhgAIYLfpKgAx2I/L4g+2oTMoWJL8C1EizJQ1KR7tX9yuc1Xx0ai/vcOnosk4283
h/5ns2+wAToz+VmLq44niglGW8EqMuJw1fy96917E25lDRDnNvmBSPwTjnHtFWBtRuBcUuI9jWkA
BFn9ddsRw8A9siM4PQQ3F2Pb+3ShQ/yY+aAPAsykx2mEzAZV5nQ5fDRt71Vhv/oXABpG0L8CVSZ6
b9MMMCQT0uxJs3P2P1NbYY+ZRJbZD2ZtAmTc1drDIINP0KusL8NOWKbNT00JZ4TOjrzWV9+fwdX0
tM/Eq25yhmPdQk4BgZdUbeE+NDBgbuG14M2tktonTP+rpq1Xf/KONUZtZQHM5UnjxbCcAX6ScvtP
JxFrId3ZIDCxCD1E7LRRScPC9WaiT2rs3E+RdjhGZli+cOUUh7PevRj7ZzNRQKxe0QsJyOHnvUXX
4u4HrdRmOUtrNExZApC9IoCyvgrzY2L6TStMfaozBt74Dli1fXdglJm11WMjegGsN3/HqMeHdI0x
SPbJkLo+XAeinB/pK6a3DexZUMXAUf6yipNOaMDIW2N2Zbj0rfkGVcCKvpt+/pqMSwsyDCvdDlER
B+izD4UyJVhIpNHqqqOR4uPjufsfCIfmXQn8cWABZzHcVj2e3DEe4NAWv1BYK00pFybqZ/bLGOOW
lCk/1H1OxLwUhPr7s67fhavDHFMSC1qyYOSWmKinafuC5LLrGXihm2eRskvBQ5Odu4cgKSidU+6E
Mx0gONj7PC8ExT1DWL5TQ2gotYng+AcVucrIbogH4y63fkctI5B86w2zMJ/7NkSsoHhAFNiHkEE2
zT1LE1GSTC7JM4FpEKcO/jYQ0/zhLUBuzztkGxucCW5XJhtbHBnkz96MbghHd0jiacK2o09c6IJa
e+FJhADas/LXDiouAh+PtO0+S6RCyIOWfH7HuwFGEWFTx0LHq+Q042wDsUIkyBTtpXpF44Uq1I/b
WfmbYcsH00ucF/XRQWmF1lMi4oj80BKtbDdm4B+lvQ34lejkoBt5+qjiIUoauwKlxI60toLnRQUM
cna6ZK+WbbW1rMEHXoAEW9MalcXdGVwKYggVW3rcrVy44CZ9etn7mLYdXQoPcXKFbRGhoSTS8Ngk
+135/RtJKG6669i52uBrb+W+wm/ZZs4qsNQhXq1LDKBZG5jtIfX/mum5UgPBmLEDDsFFDQ/FuXaX
RPrMqgcLIg3OjEv1gmt32QRHrEGSWatc/07qLSOiCY47tSkolKgNd6EgmKdzu2dUX0HoEFAXGFlD
KmUYmYjX/NokOxUm37xK0OUgYnrQ27+VZLmUCNk8EHohVG3FiBVn5Tuk/+lBAdHvkxAgQ8wI6K00
RTn86QWrrSAKTg1EuNWLerrkeC9mrZvubLXqKYJgNXz2Cm5V8J+12dnVR0onO2ylyXhMuGbNzhhH
5wzzbRprYTDF0JZH6suVqkj3oqIjDgLcgQJGHyVe/9fVFLw5Ubz92+o3gsKMbhz9RduJjyJxAXQq
xw8dsd8lLdO6eKh1d+jIL9wNlnEQKZoulmW3ZbnbW3uxwpVscN3DIISYnJgErCcQsAOjwXgrZHba
ZxrV8MnW8Y1GZIf7AICEe31cthP5PP4uRZOy9+aZbq/zc8AmU8IJPB5K/TZLMrYKTqn1CTD6GBGZ
0rODlkP0Uzaopv/TvAHkqnzV0mVqFjWF6ZeOBD271sT/ee4YxhEpRPK1SKqnBzp/LYJ3lQ4OgzHd
LHsgKqRMy/mqSIupKy5BgXP2gs1953ExgYLLALkN/MJTBtEme8NBz12JGUiJbUIu//0mMSi1O+nO
n8QwSuUl0QEmsQ42t8VdqiDbpQZLxzp9sQnm34k+TQug5P1j3Zh2VOpK13BbB/ImARGdnCZEmu+k
NI0jSkAILXHNjpHkL3qrLg1RhGotPyU6QBZG+DVfKJ/xmo+wWJmB7p3cgVL5emi0fpM9sw01qwR5
ngoOp4TPYb/ZCA1ihzGHiYmX9zx8cEhdv74815L0aHavrigUtFPwsvW3Lr0E5wW8BCkXvRYXD6sM
m7kx8WNlaJLuHAJvOsDwFIB5cFeMF6foUlpQuNnuvoaB96HDx7EM6+f3UttUbXtjX745YfuyAJfH
HAOhIYtuD7WlT3pCXjEgUq6lfuRLC4twQMXiukHp9KCZIP+sR3Fiwp9nlYFfC4HCcCKuzWKPByS7
0mZ7xgimk08LZYZ5vltU4A+FzhKw0t/H2JRpkxshmBCWszd6Ss+YhslFNcYGFS+frnjr2O8nLuWd
fFl2v1yVkz5CZ2HrIzvQiNMcLbtpd9WA4obPrhHMxMT1ED9gDNyhkJ8qTmxo+78Z9Px6v1ZSdppu
d2F+Yf7oYC0vSrARKiDv0CRCn3qxC3LTtyNuR7OCcEkIj07yJrHxRCVRFMsWsvqMG2rvvNlzIc67
F3LsvSlHMW1Ol6U/CTy69WQ+UUw18nAyAHI5oCvS+Gx5Ut/lZJgQAmgUyoNycWvutyfsTqDWnqTg
r7wKrH8JDm7GBDmK8izIqIvWSOFof/W0AVv2QGVaDkGcue7uNCw/ZAs+8OY/3kbHJi2SMtqdVn/z
mMlt6G4kCnmzondHKzv10866i3tavO14Ako18pe/LEApqloYP5b3dHnUvnOAWGOveb6HUSxemrfa
bByZ4o1RjoayM+NpozPjZ1AsDw786Swa1jbr4lFiuZO03XR46nnS816XTsPjJ5MACQFrWvmLXmP3
yFljHFcZOFOtdHamugwdNTDNDeqj5x9GZPngMyA04hJdaDWFCvGKaSY+pn0b7k3vMHQxuodGitqE
kIImzOd3CjUwS+Jx/4qLRHZm+Q5BeWg6wQujwiejVPl0ecQYrGuXc/KuYDauUXEfSFOwhRzDESgz
NnY774iU1l0U+yrarG784BHuSn413Yd089JRe6cyD70aOvuSBTs/2vzHvpSOUkk1jJYNxmmMYjCm
yquq6xewzMMrYDcm82tiGsyizTnZGRv2B/lvcWpKbvwufIDLtnUllnGqhsWMM4Hdynq8u5LXiAQL
Ep95Yh+EO+xnk1ZyBxzCgo2VLjVT+IZ7b4TIDlfhQwEtxFtJ/393Qylb/oDKlY38/EKfljSdX12n
kBNP/N/fxG0u5hr/QLxa5aXHZbaJTO+Ju7T0fQImMCEc71z+vaA6/bURzxt1e+5IeM7YJwcSifVp
YiP1FyXH9XNzGmAlXpOaRoQ6xiUB7VvOfli6v1KL9EPjSN9oV+3pbG+SLn2k0mZDEWF+ViDczOi/
+XrNdMx+bEf+h8iAls+ibUmpJVDt6KFX9XU1CT90ffg7hGF7UxeeX2PQIkZq8s/HA93g7s1d0liZ
FZvpe7bXzRAwkW1OgpNSlBd13oHoXaOWY8lrWhSWjlx7NBUW7r4C3DZIHP6JkfecEdklTjjmTkqG
zoNCHIbHE/BNFP3tMmUbeZtR3wUhPPlEaIXTSo1lBc2+y6On55T9aB79cEBErIJM/eWfT/tXbua0
efuOzCs1fi/hS8L5g9A1VVHHztVOVt4bouABSavAE88/MjWXkSZmCD6D2nu4tG8sApYaJrgyE2uB
NqyPUM/jfQSWerNipS+fFbCG21Ylf99Nlfjsop7UOB5nSYrsvgnhB+WwoQaAEAGWz8FLeQj3Z/Jo
3279wYabJzyIkumJzRcIq4dfjFHQqIn4DGuTTw9PizrL2ZUflz8//F5j8XvGjoeNaCNgCuIfhjqi
fUvqN1Lb5w2pSt9uNxgv+7UiK2e/JN09aDb617TbPvwLZJlljGGmBqjlhJEeP3hq3YhAX2htcsal
Bw3oCEAMF53bvQDpZTv3tL8XrDlAz0dn795zKUKz4GUDnF5hwTwntPbG8vb6dR+xIZ/n2gwbbX/R
/cF5gm/r0vJWgo3dJY486bFuA0wXFUk8m6v1USeqWX2eL3rVNE06YtSfKMfiGLEzgKnUca/97jmK
sh8KtZW+3JYcWZQQSW99fCykoD/GnNCaefx0s3ksq+50E46ZoZtx13vReNY1Q2vog9UUU2tG+tLo
noy8zxxH6CbT5S2VcTJfj90hGpPvHB6c8Sc2w17xtS5Qwtl591yjfuWxmCc8UvprNIRiG4mRQqdw
7I+dubT5dTJ9lT36y10jzvC/eyJJ/uELuaBfXbSbt53UzMjCLkTy4UZkihJohCwWJRnt1Abw7nk8
CbuKwK+mJbm1nMK0qzT9I64ffEkLSUDxcQI8dJ4xSBXrbFAA7QMLQlsIv0Dzpf5Dgl2nLmK6ELhv
XvOzBLfRw5X0QoqdmQ15S04zZzbiekpcYDUQWGzdvf73Z0idro2iyiUK/2/i/+YUF+tEUxJahyDb
Rzjyh4ej9X6alp72cGQ1jheiWgxeXtSetsAUxwjgEg75b879FP7abAzcDth1S+4GlhiZRetCSszJ
2BcE6962aXYv0k1zmxsngh24zNi4PWymb+DosHRTr1RX1D/X4mCG95vSVAE/zRHoGNjkU0fzBxB8
Dw/4glmzt7utS+BbwrpkP7g/nfjYEQp6kuTOXAAMw3KyMO1yAzUApg5akHfcQgaQc3fkVPgZE5uq
CsLyjl7f679/x1T8vHJFKUmXVEtcDv9H+Iwdopv6uKQAv8Ebe+1iTbVXhlA4AueTRRNK9bIF9gwO
/+jr0WTvKBG7nVk0fCLdSBZNK6lc7pr9zRvdQ/9T61UJXi/nwR5QJi9cY1voW/LACYB1D6gxgjTi
g0KB3h+gCfcpj0dshK6RIa7YYH11B7K7TRsQdLD+GclhijwrpHRXsGCVklxonSRshjx/mRQKIBz9
EiZG96QmqSLhZkFaYHdG85SHklqrfbSH8vRLhoo8GhSg/KG5bO8xIPMilGVIu/pzjTo8EufhExGX
fSf1fCqWt696eoAu6Sz0TYQ2EBW62eGgHJ1ZR2oi5je/Xt36mukbrtnFg8nzbmgGQDs/WWkLe0Mk
NAsB10dA4tpB+tX/yEANMg30UV0hgRxfo46v5ukQBtHZ5aV3i8bL6lligeZvz8pOwBZ00R2Dgk/5
A3SrHEttRZNjQbqATF0hdJ+a1L+/sJfIZgEyozdw+bUpeiaceQNLGD7hnH6Fq/57HG4N4cA3n6TA
ZRWSGAwJhwFeI8iJ4fuWZ6ckLnTaieDJ/4IxMMUhPUWSPBTEUVSkNRc/o9zmnU1SGILKp6S9DwEp
8zmL+MVl17dE/iVSM1wMp2d7JX5ydb+r5XLT7QUSkzeI3MKyoAX3SXjbX+Lt8yvjV+R/zzcv3G7k
EfOGsqf43TYXfMBEzCVH+nTy8aHN63YC4zsnx8HP9WkQQm9RnTaKCcsOq+IW3tZ6kgYzjxD+uZwk
f/5BmKBp0y0StZUUJzLqse577XVNyEWjUYQcdOzuM1QhBYHPuHGD+nnqV+73t+2cesYOAaXYDW1Y
iimTEwPy46JcTbssPJlHvg7tcS6MaQwklQdVnV0/eVeElXoSzu9qU24kzzfQ4Q2HeLJ9/r6Rymac
kDRwGoT1CMr/XxlVA1KmMX32T82ncRlF5JyKXfnvJ4vlWjVq/zIUolmLbCPUKS6hZ/s0GhVD9ruB
OBYF5OnR/FklZlzovOWExwcmFz7bXy84rx9QNeEy01GKzzZwfxV52ND7KZdlW18UKPBNhjvTpva9
DK6N0O3Kom39uzuMSjDTqmD4VtElgiHzC8HwdvFVuF+z74CljC6GwHwMdu73GRddvZYbgCbkbMx3
WE2RMhdUdtA9zdcC7R6tPQkTiWqy/M1mif+aQp+6ZZfNI9B21y9Wlo5Fc8wgiOUWCToa0PNOvZhO
dr773EkgYbnLq/5rAi/kF0E9I8l9THfONI4RPtkDA1j2BHcPRVwcddxj4PX3dmb1DRB0I8xyeWP/
L8B/zCIy0uz8oALhZMykj+TUy43phGGkDh9d4pJb3GdVQPLyz8V6xELxPpFEfcs9+523WsG3kCPb
AH6Rb60A7MVGNKkc+lUeyRwfUEVFFDDaKYXoSmJrIcJZdhr2mxyu0/RboJeNwaAzNJtggU5uO91h
go9wUv3kgRqFKFuZ/09QDyTUif925JKNHoCycFtHOU/CsAuWHA8I+9t4SJ/R5iPoh3bGWhaIMjgf
V3hdumjVeO1ceds6RyvIq6xQ8ds06KZmWfCUrBZZLPZmcqqY95tIytR1xJzcp+RFSRLnMryHQSMk
x/T3balTAzcdbOV9gyET6DMzKAbmSFLaZW93H1rLFnIFjMGd7hcHL+jx3dD8Gh4QoWVSthj1LpV4
iyfHz6JnVPu2GjUejPCZuPi5/QuMbhQcmrRUL9hyz8t05KpOCNfQhO4GYeUh843i5xrFcDsVyEJ/
6o/s5fzdqGtNiTHFPiGtxbXEbPC7VllyNzHmypGKvavKii3mswKhwvztvvlomJcluKwA6kId5vHa
yx4Nu64mSTT2/dq2NDlCzrwkMiSm5sfecSfaQ9CJR/oe8ImKJM6f6XKs8i6Y29ui6goCR3G6tHZr
8ufuvWImrR0qxVrqKV3oQSuJs1aD1drm/VDb0O584SyZW9II7ZD29jQ7w11JWZSDfsuD9jd+C9r1
LCmJfjKG2FqFb4gWqcy0Qegow39Rw5fKn8jnG1gpPM0QXddrzaAivp7BZU35jCY3Ff0ngqNBD6x2
AjOE7OLDLnwhwsA2nac+or4PWodHyk3+U5S/3GC1gMRDN23QGtrw11Ps24GiUTHSHoCsR3Xkbjar
RpkRn/V1VYrqWZnIwXxITEIpHh62oR6sq6Ccs0EOMsz4Pj6RF973DYFJlr+M65xUe13IEDkeK9bF
tDKz8Xo9y9arScgZeDSFfrw6w14eEZ3+6xJO9nEMjb/7SGtBA5uzZaW1NYP3y1B9041IrQgWPvs7
ocquFsM2M8Y/m4Bho/YbuR0AkcthxLDwANTz53Fb4IeZFOUGBURxUgQ2PYWmLHL+M08qf6Nyq8vz
pYYchW6Pr0Qbb/Z7jlPDC2C7Xu1mLM0RmSFheexCaCEvDmWNKFk+mPHAy3M2GxmkCjZk4xJVJF08
5LAzggQ1eScpW7Q0RcCxvXV8ApPa/b4MddmHroqxq+bripEXDrKAe2SdwG2f570wrtYZSy+PgJsc
bUwpgUgbeAKv+Nl6QiSL8Xxzd7QsiUxQHPwSxNTlzQea3ilU/TrEjqejA/OAtFm81CndhlE3pKMh
8g5/gaNtsATyqHffIcOlJVYjjQPe4DAlblC0cPP7kUTnvVFioaO32wK/o3d/KRAkTYvZfhtaWI4g
RK9BJETm2VAAb8GG51XjyxDbB9h/tiLziHQzSm1tTlspY3oR6u7ikzgyVXDjbCKOZdsUHpAb4xEu
qTAgy1xEEGqi4Csdw9nmbCFVrOcglyPf0B/DqhTuh30NLP6eQQAXXsx4RstrSo4QGtm5o4xkBuBi
DQeQGC2rVMrGF7TjtNgFatI2NY3Fq1r4foHR23SiBymhcU1EuKYdnNASMhpr4bAIAK+XiLE1Lsf/
7a/6iEU9FLqWbRWSwhxZ5guK8gnO2MnyTn4e/EtK5bNxnuTpZBE4n1a9lLZwiCcKBWJUklw4JJwo
NAbbpyukYpYtHME6TVsOVwkvVF6HBZngFL4wTpIjoVzsBTpdksyyr0O37QjZqsSmNrSEvyMHi7Og
sHyTUNOXUa/OapWHbcO0Q41X+aoyf3jV2nmA1mvM44vO5H97VzGlQjRB8SFmVq29oEtPWYJXfQHM
3hli0VOKEh7zrbsUNH57D1lFWbhUfQ7XMQ/F0uHd2RUfPKXPL66R6FC6/0/O0B4Uuu/5MJteY9Pn
c9HpLICCdB3YALOT1/iog/EbZScnoH/vRqzR93hroUlVftHi6Liyt6q5rhokglgmGYy9sGzvYxyL
fBx86pSgaRcbYNhyLMnWDIP9yG2BWA2CAJ2zO85fD4vIgc0fa7bZrNwtWfYq+kGVWZv0+nLC5rGO
2AHfWSbe/qWD7VXPlmnJfNZPI3Gp8mcUupKBsxILy+ja5VS+QidEtbwol2DEgYChJLrN1dKsJspi
gWuQkxmGcggcoJ3l1S0eKs8nmdSutRdywPYncGPeMwpfEMW1xVLZ8YwDUFSRwMv68Pm96RJxvbPU
KBrZ69dbhJLZ8jn1qp4Dwp9PnSEJ7bTzD3I3lVVY/ec7q0QhWARqJlb/l38lyLesjmhGkmPJNS0c
4wMXaqNaORNCpVuEibKRabFhijEXuSKe1UQ4EMai4v0gsw/6Z1jeNrkbwEjsWJEvb/40efhNi9Ol
vugfoHfeAIol9thwcDh9xEVe1HvR8XxyQWrG3pNyL8IhiF62jpowDCx5jUiLG8oBoNB96wHLxgc+
j+Q3IgPD6qdTLcoSPoOCRfjCTrAzaDZqdOAuGn2eR/FDfeBNL3lxXAMfRE1RYfSbK3qbg+dabCio
qszgKRmaM1EUFdq7n+nKoOy657q2fJIdIyO5REqxBDKKVTLe9/N5uOm5nh/KVHcOiVw7gVDPCqOU
Bq3eE0qqtiB9PZVzHezrUtmY8A5yLiCSndTsSY0D5W1TvYuUU6/rsTOZY6XJH+eyEL9rY74zCL5I
7dkaZe862+Y6hIHOmWdxhcJI/IRTIWjozaO+DfPqHV52S0CGctHHSHHli/8ySuK124sqrUPDxwmH
jzX5eYEeaa1hGaFb7E/AhLZ/nQ2bYTuZSYXWyToLU8iCeKTNAsH9F5MNShuygO2wb/jL0/y0rxn0
uBmpJIjpfcp4FymRhyDAdlyEWL+6X9YxUukS7hsjAaChv1ZkEeRAFvDN4Me64xHtxNjcwYk9SFxl
Tg3y/pKYYkBveRvg
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
ph4fbHMLdHMt9t3rD6l++tYcXEMDkmgkdD4mqYPn5Ze35RUC0m4kgOryQJwBCU+MP5iDaTYYRV5g
4SWI0DkcpQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
p3MoKO2wTFS+7WBVYUX0FOz9xBvTflfGDUU+W62MMVogCsaiuXr6A5NK3Y6MmhqxZGkElHofu+sf
FxtOG7CavHmqJtttKJfk9jzLq6DGYjvPrhDLfonBFJ7+qWzop9HKJW3IAIyPBrOX57C3hWf5T658
fwIou8Pk1CYK1P9flps=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
En2AK/Wgqk2oLRY5SjEfmbRdpDPJJgf7r2ZCEonj0CmHo3+r7CvDsdWlpsV2KlSuYhtpeX+vuwVn
2qQMzPyxnS2YcpmizlDVWOvi0zV4dRjj7r4CCVcKb/9Wg04VnnxoLgFbyxpZ6n8uA0eWuwHzC8Yl
Z8dzu6JMOi6EO/x4ZcIiI8MJiyOboyVzyx7V+ja+eS87qowm7tAroCckmNEYOvARBFQmT1AtIHSy
dyOlUEbZIpp0vqV6OpKK6Rr8wiLfCKJqkomGF40yx5rsJ+8bNlgg6udeFS0x41q6T3//RHoERzWI
FTeKY1UlAiB+ytKEUUtCnwQD1iwFGQgfJ0h2Kw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
fPd069tEZZz5v2NgXzRiuqS2lAEPLCdDDXFukVTw71UsqqbYLfeXFaPaXoa02TcQZrydmutcrtlR
J/26u3DYVea+zJKTBjcHqbaopWcTiU18NJgULOCQOWFJqPgyEhxXpIvd2ETbgpM+ifWoInP8dUlD
8GhUSqmk3Zup15GmhfmNSPFeHlAaXNEYCxS64VLPPqO270tzzX2ffgkpfjih3XEBOEWV2/fRMEIU
3Np97+pUw2m+IJwt/HQ4PJVtGygekdul8yF751pcjPuaryGDM85zzRgGFhGSovp6sBFcDSlu3Jvt
adzhldYd0ezTTk4relN5Br4pkujkM6OY4X90wg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
tR7PxLcMjSI9wwUgk9tTHdcY8Uwia2NXW5kaLvO9gswxN1GtL9GSPgbb5zr+sTnp/S+LKTI+02KI
TMB2geQgK1pZkvdk0+Ol3vq6Tk3Zk42Qe74Vf2ZvuojvmkV2QKZFg/aa2tb5O17kne5a1IXrg8l5
z6Yi8tPHSXCNwciJWpk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Bds0en+2c8yztwhHVpMedOFRj8NmE/EEWnfaOlQDyHm80o1CcC4cZHg54ZpJfMa9/U+YW6bNpsqS
FhcQ+qEiE6QQJpUFJJDqKhpO5QotCv5d1x0qrjaitJ2226PAPA9tN8Z/ZVce7wJ2S3dwf9yv+8dO
rbJQQd2+lF8shy5foQRER8hcOnAeL0MibzMiJVU86M0mN3Iy0EBiQ53foAu5et5iMNly+0Z9/L1h
C7LP+1MRwZ+VA/mHmo+cKOnpQvLRRhGLaMCOfV7WF96dPXwZ3Z0TmQJx7RSddqeV9LftOvrNpRPm
aZmc0GNJbK+RYV604McyE2SwMEOkx3LMghALCg==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
alO/bSTeEnbogP4KcCzgjgW1pQWnX9Bgzz3D9ibL100OPGDpXUyCgBBmGhN1F+GR4iwTbtF8aSP6
YKMJKr+0QUueXQWwattLlV/7yK4r+c6cmCm0MCVhnSiJHVen61GwWEUTqOKfd994wP7ZJbNdNk5n
0JP5kG6akdfavqt2saV1wC9SH3QphpL2qBB5dgec2Wn9Z6tERWnKrNCXCbntKuofu8/rom6f7/AW
I8Dd6ms+fvD2PL25Z6FKZSFzf/u0leeiQUpvB2Mhe5gCIymdEICsjronnhzSfBZmmx1qDmPXHc7L
uU6kVDl3MNUB3mCc4AvJCIdEErJ1cH9EPBaf0g==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KCBkW2omby+FZy53+sB2qtEp1Oa8tM9yMQWpQaEh4yvplMjPiDdlXmiSm4hbpZLfNX3IaW8TSza0
oFxVjuH7/T+WzbOgY/r6i1SoZuE8NtexB7fAymGCfsDcRvuRFBDUt9jmkNxiuuHL4aVNl5gU67Jp
sBl16ERKxQGL94PtR3xNLEYFXxkSYXrIciqnbXyU9KqS0axlAHXIEOK7mm/hsRsRj06sh0uSf7AO
DH002lKncjh5xlS+ad/B3fX+vaA1r0RdEf4gN1nATKsquH+Ezcunc13CjIsU6WmSMjDcr2wjM1+V
x5raLGvn37SSxXKBZRGMYMEnl+M0CNQMgcbI8A==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OKpvCZ5EyJbwgo77eKHb/YSI/lADZw0WqLSeEIH3GOBl5NeXzWp8RRMTLyWMYeG4JehSE9jn1nM8
FPbheCZKwZBAFYyZ4rgE8YGf/ykvuflSJm2uXugw2Cn/Zr84QaKZ1e+OCPoqJXO7IVVpzu/1/c5e
t199mzUJEQbmVnBy09AgqYRqBFElANrfIvkBxa5u2kh6Q3gKrFXeXiFGDdDoW9xvShdZClFR0eSg
MDl3FGGLguyTSZWrFdkpgryN6kpruoRCKFntoicEsRcte8ecJZhgcNsC2XMgZHGFHn4i+mQSQkM+
f05kNS9z3oa05gupkS5T7eunOYwPfeAooMVZHQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55296)
`pragma protect data_block
RfYxomztYJaIWoKVoB+VWjfJVcP0SVl/YWtolsE3g7k0s10G3jNSTbPo/Iv9J+PV/N+HJKbDVzdu
UeXyV0zXlVw0cbtFJB3HpKf1A3srjGoX/fco9l1Q1dfXDAkFQbkm8O20vqCy4TdvqxZvScC+UU1y
p8TNf2DHsvHYfrZxxXtmcAcRmmrW9EhOjPLXiabWoMwniXEQjzmH3m76cV58IPsCi+yKqjDQWtN4
OG00VnvmouoKwKOAxjq7OVU3yvultvc5hJr5YKhbW1nZlBA/7jdhRiq9Lc54arUxWoPfHhJSibq8
J7vTHN43MoiN/6QrrgJ74rd3+Qdm7U3iaOEmMu8wIOEtSlFhGAV7ZwHP2gOX6Sh8bMNQLLvv8BbN
J+0PBVH5abBt+wx8uI1/IZgRUHrDO2OjT2QPgRyQ1hzI63VhC3SAlDaoC78jOFZgc5if0SbLPnT3
yD019dt0Ycxg7XTapAzhg1BlL45SZpsMSXhYK9JwA1ZZhQRallZUe6u5jPDPH2yxtPgpeJfrSfGQ
oP7w1TCb+wfHog18jC1KWeS9/iclJEnVghZNGowbBS+ZAaaJ2pQlMmjQfjRpzGBUhyZJnMKMWmHa
aIB87R/8XzV8q5MgIjbAYdTGIaNuSBxHjudPcj898qBNEo67mo4AVFXXIgNdRxyBTH5UCOC99CPy
LM/vJeWDbwJ0BajjxdLO5mahhS/L6OdHGlGXj0E1fiILhWbmm/IB+cZWsYEWoNFgaXTvSfcEqfcW
gjdfQFmWYIK6h5I3v/DvCbPw0ZWbQzylEG9AsqdBmQBiRYGn60XhlZ5Zx09wUOBbCji4Pk0GUO+M
fHUJs6c1aDBEFihGufXJ7d+vh56RPl88gJYeWpLpAU0pPAnVWOvnddDYXgRh0VRePsto+1zJtVvE
tmzaI83a16xuKYOQmOySZuo3ie9WNCPrGBCTZ0xRnaKmbz7B2a2opPANit4CGIkz9dFECfx85hJg
TaFpTxOZE3UtwxC8mb/TJvZ9cbAT7DuEb11kREXS/zDBAKczHPyaDmpUnCQb+4XK8WrtumzU63pJ
YVafSAqClYVHio5ax1MhKLBOWUYNq/PpBZn0W0kUikIOxIlNaklvbgZregyripcOSGTjZpYsihNH
87Ao2Mbok0a1NJWfp0xTqSfhTXH3sGM03tIESEFUGs5gVS/6oFAAe6VXUAjdsq2tgGjljIGwGZCC
nZbzo/PrWa20XaTKFJXylofwHyWXeKH6v/AiA557husWphy4GNqsNEGPVvLS3+X+PDyAp086njl4
cqoFJ4xbnwjkzbjGH8MZB6d5xRrf8I4PtIHj078IQM7NyzHR8S9IhyL9nTxg7kFR2ZYL/Ex2D56T
737FkA3Fk0Eept3kVpfDawFUtWXEMa0oIcrj5L1qn83GoI/aHvPEj8L2ikRp3CzZlF9OmLqIDzKi
AsGouThxQBBnRrdDkMLJBqE8SbXtQ3cqV1xkhgyolRGbmz3yAUVlgiXm8DUH0JqIg2lfgVI7SJ+W
rPmgKDLGchFcOx9a5W5dU3GL8xnYkBIkz2fQ1j4UkaIzc/edEbqZMH53zRW7X7xI9TMbAywii5dK
bkzfdGoDSws0tTsA7Xlw0HYQ0+2EeGA1PyVWFnmnHxJroZk+PCrFVjEqRxec5BPxoo9LcT8ahB2Q
9zRihKoCKRFAWpA9jKtGcrFo2CQhCLJZtPtFN4pTyWx9EF91P6WauA6sbnN/7rgUxgsVxUgIT0Wj
aLOZwTPhc/5wU9MnorUHKGVYXAO7EvxR5j1MyblnkPd51cjDrHQPa5tYmAeUGWxoAZ82NhdY3038
S5ypDQtPFQExB1gVPqjSZGJklhcOdlCKDbWYsK96aaB1Yrwp7MoYUKn2nKMoWNnyTGgpYW4U7EAO
GhMSmr0oUk0pNJzPGp7F4CvB8WljOM+Z73Zupkn4WKQ/NVm3oULZYe604udrdVOIboYxls/5D6Ai
iYmftPkqXM0zMR1UhGYbYLps5jLtgYvlJA4CYjizVQEjsQIJQdL34c9VImSe3Im7fQQkWxJ5Z5WO
3fDqfh/a3yJKjbbKVJfwPB2R6UV8fcBtF5ks7Vls8A3QO7aCMrT3k84J3sKuhGZIegLuy+DFSSAm
DN7dKjzeYRW/mk7G7ELwfykbUmKnN3C1AbfYPi7fNR2d+59J2/YdZnjEKjlT0X1JnWZMIxag+BzK
HA2+U3KGVZNWwqIoybGhYRuuXSRhtgYRr+5Ix74XSQmO9ySH+Bj3pU1xn8BQ8s0ZhcfCHBAGyASj
YgMajayaoea5paPsAZ/3/kmF84ftDCLvWY77pKAaWcgroVSxWsUvdG837hHuFRRYbg/Xepke1S6y
YDwA0UAKHoZCHpb/SU6pZU9g5HOfet/PmbtX/VLWi6zeBNtgbh+fgNAbL9dpuztrH+jO2MWHXkMC
sNkX6Ws6tZXuvFQIcE0feZ1i5neMbuzVYql1T8Nk8jM4oV8Fml1tX1ZucKkfd59nyqYmlt4pCR43
mFbDu4e5Kw07HPc3UGzO0TvK6005T5fAFR0kjLaTmfEGyZJXh04rk4dt6QjBhLtd51eF4wYjZNVy
HYMbZisQ58Q/3ej6k8ll4vsySbbTggDyKw7D23jRzz1Zc3Q0CjAzpACgpZ9LzF5ryQQWqavR6xyO
xZ6bGyeHdi7iUDdf85z5Q5jlFSGMD1LqoZexGKT9v5HDKgKTxlfwQ5vMCfB8AEfF1ABhDu8LAdcT
/TZbmY4DmjLlD+jHZdLGkyTSgnCYQ08YToWGbaQ876GSHOtGOud40lJHfU7BKQvzmMlc32FduAWH
l68DgtICMLFSy9vnIJ5+F+RKINkuVXkr1AQCr60KA9/hHF8iobVfaoFWJFz2f4SlIp+MivqX+Hhr
0Hpbq6//o3L99oiBzcdSSMYS2VCBhN5ubCHuNgV6WYxmx/hwQiWPBVu+AWtqa69/EUEw+X6mFoKc
QGiHC/MOQ4YOIMQVgkk9JiJWgnmxGmd0lyiUx9Jp3e7JfOE1vk/DdemGzdGnIcXolOKJ8h6xTFPa
F8XMjAQ56iSZ947nbQPjaavZaZ49LXXySNZePvmj7aVjwXm+h3e48QzEhPltpP73WNCgyrrd4Jh6
cKuGboWE8CVYlVezaGN8b/pQMmvQl75bXvmqjmRucR1N5SPHL91IvndW0IS5mirUwifmUbOGEVXN
Kz3F1wfyrF/jFW2ldjmHL4GP+wVfGg9i4DNxPVzy31eegvPUz67iCUxinFvClAnK+5I5vynb3T9k
YRyf9bq82J3AosKPfuWe83xLaSiFUFEcv8xIukKwmK8jRqwmw/w9gdcKbwXvmKtaSy5D5bbsg4Oc
wXkFznkqDFV86GxVXpaNTZNrceWH7fUYTmp7c5K2c2J3ClemmjoC2gEFY5K0USbGHQwcbw3tSU7b
0HRSqdriHISwh8gVYeB4EVj6kWobVa2wT6i/aOKlgv5geySQ6S0j9KqMKkeWG8PjiIb5ytmWIXsE
jDlJ+m6BN/10j9l4N2hZ9freScshZQC+8cdQA3p+wo1q70CetaLeB4EPp0K39ct9ZxnaHJYjWszm
WmdRfHHuLPPdAVCe4ql95qEH/e4+I8JThjwRM4d3eIO993Djc6KOC9Q4JXcXKo77w2JceK7YQcNM
TUcbJrjw1m8TsL22P2Om5oE6QXN9weqEr7G4ATg4zjaFqcDlPLFNvhXS3KyTpP0mBIrWc0mc10No
xlYzU2SKmXJ0dlOBslw7gMI2O4q0bxBosC0NluiY2o6RyN4v6/8Vy2HNpaQt8p8q7lNE3EONtqgM
HwmQtVa2MZL7689je9SPUEgpwI2UsoRyMLEwYjmB4vGsqjM3sFfr8+C5Dvu7BN0CDGLKwCAteP4i
ZbDbA0sCL+rBdyTyZsrHFJPh4+lWTiwOwZc3rnkgQOwJpYY2bFj9GpCfVJWxkKs4sZug2PfYVhSG
uCoFzPKbIV5daynqslfES4qq8VQUO4n4AZuuIPBkjNNg5o4P5VUEPKCCZH1crektnsZCcTHuk0IW
efpKmZBVI7l23BU+Pw746q3z1IyMWLy+wJl9Jtxk3y0iYWjLrMUyn2qGQ2l8xnRhaNi2rXxEPH9Z
Fdcgx2+9NQXyEOyu6OfidJAU1/629qLcN3vxBCAN55RhY/9hKMo7aCjeaRZAz4/C8DynVt47sr9C
JkCFOqSnEsn+2soDa7hHz2bd187BmVNmqaRWiiJrrTNksuHAh+OJjNMJKN4JRNF2aB9Zf1GKu3mv
qlBoFaoXisNyU1JhY/HOP/OysRPLicIgaHuCjSllRn3Yy7l1YWMZSEMOhAtIgAjucXO8ugMK/+HF
p9eFepVtLCnEbZZXmXWNg1TfXxWebPFezh4jRFUhta3dTRcd8fe6yrzrTwOr/iarIp9ZeThXnVMv
/ZwZUN295rmwWOQSGLTvdsTkhqaa1L9FM1TC496BGooao6a/Ahb7N4FrNVIJTiBlLz5VMWAipNP2
PwkP0UU/VK/EVIwF79CnR9Yrk5WnOvVtQQnAuq3Aw/GWCyeDGFr9QhiKHVCGrTDiv0Fq8TNTxCoA
TXVAtX7cod1c6KwCOf+PgH8+sOibHs+/SWKn60sOk3Ffz/oVQ+vDKmWwRwWVkdILAQxouAS9eUch
EkJ1+xtsF6juevVEL3+/oorvL5alkNBvDlrgfhy3SubBfttRAesGQHXs1DQ+Gh2nkAVc5ApuDbwB
9A5WrJHixbWT0XUc+DEQTIoJq8V2LHi0EuhSeMt/b3MzO7Tf/fiV5SYde0L9juhvJpFyHt8gp25l
iHyo3QxxnELe80hnlARTirgQ+IHI+Lx7k52XxG1BAdK2kJjtRbxSvrj/MjA7mf2KNhqCL06TfMHn
eRKBbUZdxyDimXS14YmJ6wxcIXNCAaN0isg1WscFIo9oQmiDt/AE89BeGkpZPrkGEI3X009egyDu
3Qm+ef40DkvKchDVAmjtVUcBL6mXYcObXSE7M+unOgSln2oJAEQJH84pHZx5skD4UalkhhWCFlCY
Fj6PZSWqXLn1tIjAYYhaxiMax+P9LikdKCsf8NOleoJiSeeVq2thhKP3QkAJD/OFmMMxD3CrOzrI
Vgqu4pjLBh4KZnO1FsltCMTyKuYTX+4GW3RgTiyn933bK9Wfuj+jDOqAf7uW0GFTNdizFvcNZBzr
nYhXTzWuONBjGnh9HUJ7zTCKFmlwKedXKaVNxuGwDMbbIzLyRiElXOjFzaMsYr8Fu01e/v5hVOC1
X7nsC6g9gXRKlhYhuwXJMupm9CGezlfX1KFVP3/9P/i3pJItIbxZK2tL6PFE8KX1qrFxpytyRYWQ
mFyq24FC3ArRLPyM9ljT3xPkMEVN4zf7+r8uSoHucpMmAjTKVdN+KgHjX62n60HFTrd/AOQ+eRsY
X+m6wgbhAIGjGyYgb9ycocVzcenlFFoFi2jyVhnfTkPFI7IffBaqpyH+eJce2oqgXFBXcAbg+d/M
lapfoNws5tv9aSs7DNW2Q9pjXR/t2do/iXA3aAhUJFbFRQVO2vs2ZB6whX5qjCe9lTu9HuWS8cVZ
zoXne9g1v/eCSxfYg/POOfnJYSvi3lUbEJo1uNoIS6MN+lZpEdOw2SGVYQmlUg65w3bKZDRHdt/1
hqq73z0LCkMn4fW9hGMnEW09OI4BFCH9PwY1MK9lyxLwmwGhDdVN70zBNp3O5fSmsgjCKuXuSm3Z
KV7Cuos+9x5Ok73s/bRQ+pqqYfKy434D6ZhjZpmuXov/aCD387bgdssW+FOvddMic4KOvnSAcIy1
Td0hgXztY333cdGsOml+lCBE0vleTayha7zOAzoQSEyRwKBzPI1SExPodaMhS9637LLYtYYHuoae
DVa87Meit9ZYylH7rxcnNJzWL0JN020qiNXV5MSthJCCc9xcA9c1QjexxyCHgHrt+Bm0t8aMs+e8
kkZTT4uarWjnZZ/pKV7ehoAe4hxKxqn8nF0vEXdohUgXwoj7Yc5bcKN/3nvi+MT3lotjxHcChcdb
u5H9T8EdTSIVfGEea2X6dY+mqEo4K2/XMFSS1W7tOZwgPN12EQpb4L+KJOatoSPbTgCYJVLqQ6bG
SLy0xG9LVM1PZ/YbD/e/RI6OI6vJxXg0RL0I6FzVWpBrdOcn81mGTWxNSn1aa27dZ0y26pe+MD+C
5U3jVL2F1dMKtdDFGfSacmPDFAOOqeB8tB0U6TZW8l6+7XeBpVDZDUx9HX/b6LjqYc5jqEHIHo9J
8P5p+GbfxLTfHaGg2oxs6D5ypz810sVnG4BLQNU97ucLvg+PHWe+Z9zTFWE/3+2qxHoxOM88WT/5
IpaJumuS1gesKvj3b1dS13VW57PVMiRZrz9WvQ0NJjQvYTe22s8cTtufZ3mgJ6o7jti2f66pnJit
vj0eOjmVz9GGzOpGtVH11s9VTIU/bHTflPaoWiLZmQ3/ygtSNEASQFZFQ8JXRBPtozkjCLrGLLlv
QCyav8Qv1BsIP9fJA6ekbVOuNwk3k+Z22KTDuBNofYzkFUKR1qU/ZzvPJ4XhsTcxxLrrxoyy1yh/
6ku0pQCXl1G36LNoYj9tCGlI/A/i9eqb2o/F/VsQYqvSVKcPuy7l46pFzM/+fB2qA8pgaNPwaS9D
5WhnSg5KxVUVipEHU2+d+NXFeb/f+iTU2FW37jnF3gON9iqnpnzodpEgSBW8VChEVuYFMQSrdcHY
FPOT5/OAoo2cxoNrCap2MJx3hGBdrWDrXDTnHF0UFn2zJhqc6RfvG+qIUHOt1BVig+OUhP5BgRHm
Zw8VACMFKLwno/CccLjEIzDsMDG0P6ZUCMsuHCpW77MyC+cTAI7jRrcB+V8+f6z+KwlF1V1UA7ad
lAmCbflx6B8vPn1KYKTym04r1RS4c0uqIc+dYiM+bIH1jMlBN1qcmMLmUaiBCVbOG1I13Dgxm8XX
pN3vrsWONIv8buepXbc14QEs9wbo7zlKwRTPDsUyzm06Da1p2MpTG3c2vEL4jyL/q2CnL0+bnxTu
LFjDdMIWA1OY7sVcrm1OHzZxzrQdZoxfz9vyKdgHOlbv2zGp+/h4h0y3MStz5rk2EBfljv3ID6pH
sUT98SovdZL7geDdfbJ0zeY0oX/HMtDjLvo2eRUGjP6xbaknS7YbgV6GWkYpt3rr3Iq02/FJFzM/
zBHKAOJTPPURqDzdGIxRapu3MSPSksj/UG7Gxw2oATUPYjFjwS6FBk/KM71RlGhtTC9aCIEG+vrl
+OhhALwqYx/xxfI9KEjYfNWcKZu4LZX+8eF2lkrUqGjLhvPYQmgxG7rYcL3GHsNS+/b9A5WqIteS
19M7V+bEn9oIHn0RDZrbnhNPMIKsEUoXLSuPmNC3kkK5PySkUEccWghn7nnwfKhp/4f2nOtIKHjj
HGDk19v6ZNxHDhf+bBlKW6iYFSZmt/o+5Z+7NiN09wcBeq8wcVDURSbnK3PL3e5p5EjCZRUdPJ+4
otfCi4csWbbiYPdFV3SGAMJ4n6169uVVlEPvaHJWam+43Vpm1vvhikYWHtRgZV49osggbWGG3m9t
halZWnsOSxuzt0s9JZs9y1eq/cqvICZ5FeR90JztNxhjITxQjYApc/0OHLd289qhfX6pA1PTMIxe
EjOKhNIkfBy5rzfLT9mJhPjU/+aEDeuWYpGXYk1zott4qZEVRez5ZTwK65822AYOXXuc6rGEmdyS
MVxin8icnDe3DsUBvuwhmeILrJJxTXpGx/wflNij1vX9uvRLLO+tAn6OlXwtRR3+mV0bZaNSwyyk
oRe8XUbovHjN16Y5p6rqZ3XWU9FFRKSGS+zWZQ7U1el6X9RI4cfA4xfNE/5GmQr+GZdkXVG3P1PJ
qM+Xli2S8qcKplI+JkaOqXmE/4532l33viawwHwCCbV/eEoqyiFQYZZRDoijBQbhC0QfV0n/kjDc
tQrDhClV2mC/hKFdao9PU2tflj50kmJgZBcs4q/OMpvNyjKDE++4Dk68ncYzxqVJq3n7xrsdXBY8
KjA1ZnrdoA+nxMX5jqATinHivqMW8Wag3tvlFPAu4nLwUhZUBmH/0Hwgwf2yJzIvBq+kYCpjOOfW
qg09e22V7/PYqFbrmwaIdRy0BIu4eR79RAfNAoLbakZzyMzdXBjHCZQcGoiqCO+AqbqX8v/d3qHq
eFYaY1ynmwU4agMsIasdAH0BABetWNXsm8IL3oslbvIQshbC5Vx9qcgykKJt6LFDs+9o4lczpQCV
jxWUDV89yJKWgechLe1xh2A2s32V4FA58bpu4NhJVAlWbJ+VFO7JFcHJx1yObJeOrnUVVJJUUCgY
mciqiCWXda78BbsoiZR4rH9RJDZF9dGDBbCCmkaCTELhnQm3cwEXX5PtXl/S4Q44UMn5cVJIjsV+
8tSACs7x+PiIBPyyG6LvYj6Y2uLFXI24pT5KmjO8eT6AsCzBMW2UDJy1cHU29/ufJoTCk7O3lN0k
4KPRmFte3VrnsRYQYO2jdc90LoqtidSQobxt9eDzzE09NmXk8Tz0QKAuAF1bCkQhB5ESdAtp4U3U
Xjwn3RXzDkBXe4UE+vJRLIv1p8fnho1oDQL+AfdiisyI862+XHwYK+BPwOyXAchUxBq9Zk7V7V3T
Jhh5fA4nNbbENi9x4epoo/7CP3JgjGq1bnBFFeA+eZ9rwak+/h9OOSwyXrp9pJCGxdYB7zSi3B1D
yoPkD2i9EOgjgAcAn9Qil4YP5dtS91KeioQQz87/c9qhhicrrxPUHH77f0QuqXFpq5cJi5r0ZxPk
YmLTx2WTVU0U7toQHmzYpf8StySqDIKJRh13dhT/2OGHs0IkGBGH5Wsf+PPa7AFG/Df5xkaBULew
9UKe1QwEvtXCTaaXy4NBg75Uh0EUulDPIPIB7dAuoSGwn+iqHFUkdC0PF6fPq5gfolZfsZGMt7kx
QZdOGoc/No3MSQ3ZjNHVr+nz6NK5T8lCFPnYsA3hmpYhk+h7Yt8N4DB2AOfWvl/VpI6IyYxVd+YK
ThpO6sVyn2ewQA1CCkqTz4l5t6v5x5qKM9ELs1s6ObUvmrMd0kxhNbaQOQvF4xSM0tCz12XybaF3
MVhJ0s1PYGad99l2Zcu3dwfwcAgfWQ40Q8eQWpgEB8wt1sqkq7U4oxRWSBd9MvQ3zQpV8xkOaNxb
iosKK0mLGNbn8pOqSH34gPr/Wqt8RmFNcOebSZkCcUjQhU9b2bQaDb6V/iX0dx91V+TpMmsUPj42
z94j8syU+gJpgewXGBI0FvJISNxosFfgoyQ3n6mncoLjxP2CWmTZVHP4BbKFRSkms4W0ZES4mk7E
aHXzM9vHHETc+yNUaTNmdAIV59DxEyryEIvF9gfDxHTYODyB91W5BeR0O3RKfUk6n+NGZLoVtvgc
Ra3e8Nek/Pbq5kN4sErvsZ+QMg/DLifYf5BQ0/4oM0whTAOxcE/a8VmYnE5rjPaevw3cGK4LMvY6
TN+HZr2xlHm/Ke2jIVI39bz1oo9TfoNN/fsFJ4Rww4Joq6/k/hUU0+8ee6hVWGs+O/CruNIEIyRS
ckoVaVoUTkIcxAeTwGjD3+HFW8e5JTEf/1Lgyx7qvplyB4qlbrqVGvY9ZeHZut8Hw2LjJr29EaOH
eJN2Ktioh76pBjYdQm4Ft6Hoo8IDNgkDsuIDLUCVi5LmzBXNJghq5IPXcl9fzvGJovaWN/98yjb5
Rfkdqfu3N7Afa2E1Kxrg0ZDMfghXLYuAn56SN9fcVTQjtSEtRi0ha55Und+1hODjjA/Bbp3YXoo4
9CbNVnOHTHuzTrR8zwNuw9tOwUA+zTV+yR8jvEj/80pv74hKvPavbakA+kbk6WFQxEzdU5pbeXaB
SR3ZqOceb8Lu69XIxdOCNvA9MNRmaBBxzYCc/SvRC8uwSdmUiXvAX/8pnWT3VppzrPIOp6Yps1wB
tCx8dCUnJht8Ar23PKQ7qpRQKKfMOH5Uas0i9SZ4hAwqM32G5fpO/w4QYxulbolJ/3E5761Rtwt3
rKB66C3SO6i64H+CAgU6tl/Dy8sxzvfRix2JQyeRRQGG/0ZBuwg0RhQC9fhMhOvV5CxMOrKTDQYN
kmKhM3QToqET8ddWmRqLSH6HLgV2gXg+kr+e3NTf9+7Jb4cQbpbufsO5wfSRfvTdCa1GmIo59pB1
b5OYDqo7gSbnShvMTNXSgY+o9ejChdwW4ZD0E0+U9OZ5SBk44UBV4mqMmcwkWNA8IR8vIW8pOCP5
0Qjqm4BSlsexA0Gr7/xrWw3oVc+xa0EVW7fBaHkcphyqMlI6Na+GqqPJH7flSF9fmybvOEbp/6iu
x+/j0MXILLibUY9A4YotjGVzSlgLTWpE1U3x2VX++k4F2/+ND7LrrRVg4A5B65TQsXv6jbh56QnG
mxpEPeIITwjlJYajpwcGi8eEyEAHcylOTUoOetzMjzowEh8gYuiGNCkOOWGLXoqnhoZjt9eNxtaC
4aJKtAwYmgmkSjb2DdGygFSXUI78S+iftkAx6nz9yKK6kuXZ7Teuv6Hja/qtcGeSPMa50yHrx+v0
cCG4a80NazlHkDnp+FyyBj4kZlt1kFcvMRLGek4KXGKmX32TDn2hTWBO/eI6VDNyPasW/JgR2Oen
hxeTDzhNAOEkfg5l3IOeprwMUtN5QIOcyKV2ZzxHdOVHOVV7Gj6DzKklXGBE7JEYYrxmQzz2w3Bl
bCKf4Epc6AadbrcrrKNhRr+tOm6EsOlsO5VJabIMSTsYQm67tgXTs6aq95u5CRWOl6WqDeFS4jzt
4SmMMf1Eq3sdiHQbqS+7At86FYpRTqjQhqtn82q4tLyQiansq4m9FEROquNDX5kk9iJPX+xjGQ6r
JVbwynaOT46AvXQJurdJNYMwSPSmP1t8x47F2Df08W95uOyEA29vx7ed1OqBXBBEQL9TIeS55Sb1
wOjmSh8JMY+wyZc0i9xKGZvpsX58CMBASjzrQaKb4wFvPdp+HYFFACqpzrbQ5MwNJvtkhfXn0Yjf
vxE90mR/tlCaTurMxEOD/P9Uq7PQpKVLwrOY6U/qBOz5AhJR4w9T73MztGVXIlTpnGZ92kEuv/Ql
ZCHEWLBFU4ZyXl7NedeGKwI+py21FyXkWb5q+z1MOsB5Zmva2gwW1q/4x0rWIlHnF4dSpcVsn0OP
SFirR/12DadBsmSOiduP1lJ39kMCFG1g/5MFO4pl8NExS/sietyS+QMaLeESaGEU5uvt9Gz1bs9i
Cl3EF2SkVz/SzsWlERVhEhKyBiJqbNdEvRBzkyrtS3CBANV65vUloOhaZCDuVT6dQ8L8cclgFa7m
AU2v+uBJ2GdmR4AmzkoXmug8T22sHDSjR4/asEn7E2LTtijqLNAJjx5SvgU7282u36EtZgyvxt9p
oET8SCQaLXuC3nNm3lkWq68hrb4LVHPiFXDV2ynegJNBfQCwDR7lkg4+hpskepIoDu2XN8COTwVv
NrKBigjKR/sDOnZDGrMsFb0bMmgg0WfEqx0+xt5nXp5eQsMzFnmvXIOQGM4T+DEkKwFD2CEF9hpt
DWhwko4XAqXAdwi20tOD/iK6XUGHlZqw6o3w1PlM7vG5pEfEpBvlnSycQmZVCYqvR7gL9dBz5CVw
plaI3MjkruKASPIPy9GmcznfZTJZ1zruYaT+ChLy0mtEpq1O1FzfPpvXp7Nxn5kodZ9gHnPvYeoh
av7Z824+gcNwOJ/kzjVi9inlSvF70pvebSph7UFhF2bdfvehRlavnNzQEx237Ov5nd7VW10L2HS6
X0seT9CTxcszJRjRTvNjVoZDLFuHGfCVAKk1OgPoccCTmgTy0cNs/zyAVnNQ5xicbESd2v8rU1HI
1ADG1yh/ch6osHLLo34JGl1vnJwiyEDoYy5k8jk3s8xAv6msYxbyOn9S0ARvrsJ4JzPnCtpmezFS
a/r7vEx7Yt8bmJRVMTT6C6Ahxd2dmJqKNLltNPed96nyGhGDKxLpccgC3KUF8otmJ9PKSPBt9DRj
abig94jYHQz7wl6y/3ss5UOtxve2vSe75bXvmCHJGTxq7RBvZPA3bn5FEJqzsmkO2SZGQ3GvNjma
+6cQSltREIRvTNJSoVbdT8hDAE8GM7JoYZS9BbzgmSWJIE0UX2fp3pPsTjee5rwlFRgAvRLUI+ys
3UwyP5LiEDyZFCWSasYIdX00VfGtH8jT83GSO7Ilb7jqp6dFgwh4vFxtrDI9CfAndO0ihb+pEJP8
P4Hq61az6A+nh09D0z0m/i/Vs1XkMobDMaHzpjizFrUop7GVM2pLhkqsUmwnmRDSeWqByeiRVMRI
yGCHYvK1vOkP09l8k7Ct44NaEg9Lgz5SL5Dcb96A4X/+HUGbSVYuHh/4WJtntC6UW5TStqR7wbxV
LJba4NZS7U0XPFkPi+XT8SVT6E55O+Jfof2BcwEXwIx3EwlJ4Z3BcyI7nCqcKPq1XaGAyBDzDhzu
HfbW1fgzwt9l9ytQDD3ldSMNeXByVkVwAXnIJlJ1zF8NKpUTKVxHVE8iB2jVMAukFvX8LsyOf8QL
yQbGuwJ7FeRmaukkBuBLUyvCaEE4s+OmLQWD6gE8e4CytctnWAio3b+BgV9F0Ie5PW0WidHCdssF
Aul4YDRecDrsNh5lgmXVUqlPokSxe68fSJ4DxYrnrOam5GJq/bmNC+wAwO4R8IWC1d4/KwWvP5xG
3tj+I67D0YQ7o25zvsose5owO//pvbfwinuDNpmhqK59o+vbAJVwZEwB9feF3VzR15sKMsGSvCxy
k1sAIYh5EWSQdv85hHgKOO/XwbVZlWvdnYoSYqIUeXjt0N+AJg0TwDeCvGcQoW+aK3c7kqY/t9vF
uAC+8NqlgSR+9FxBFCbwv6Yma/CInqk7UBA6/BjG5q88DVjnt7wYRK+KHGdo+KVcgYC44wVDZ5l+
veJP/oQ+02WpnR0RQ2giafiWaGIWNYxVgiUM0XlCT2CD+ScQVtURmGd9o31RiN/Q5kdejAn4wRWy
AYqPecN5wxQXzdMGExYBCmcfz1b4Aid9w5ELTpX7/lttk2/xXvIVBrFuVcw/4BQY2GvIq33PiQde
WsCYcmHlfJ8zSD+fq2AYwTLjtHGo4Dw17zPQj9QR3wPWLPmkz7+zyXEH65n8fpQrlect+aR116Rt
zyPLjzcjnq5tDV+fLcOYephJiDKwriToA4Zkk9lGItLvrvNDWbqBEnjaXAjctdhtJ5zLlDnTFQMI
dpiH9Mfov73/z0RvP0O+YstRlkA15jr1c99vwMY7Mj/BuD1cx6YwclE9Vr30Z8M/4qGeBM7pxB4N
Y2qjCeGkka2oYC89SQ9hBIgKqyLraClWjIi7WHoJOEp6+9id2/rn6bnQoN3UrBg1igB7o5O/UvBg
ntqpODZXMPSEhWOOlUCArvEg+mYjTpu8kbT+Kjz9RDwfsN/0RHEolb43OqaVP/kKpubNHoa+45Cv
oNLFBJWjOVjk7lNnVxIKNK1PlQtbih1faHdy6QkpqJSFX2AAM0cM5ndHIknCpkp9r6Y0nfmh14lF
rzzi5VOaHSodR6IEThCzydgcUspsgeFU8+5MtH62N2k+oQrcn0ONl//hKP6rF8XITfzP4xs2EVJX
g5in396X8qgYac+HopAkBTe9fPbsyjJaVHHw+wT2BrP5gVsAmMP0nhWDMKP+t6nxOxJpH0pEKeN1
tz3lsnrQmHsnk7pRVdGp582H2cg/OyDPQj0RarUNHimqsBc+Gxx5jeHaWbMBXyMEwkAtxWKuW5kA
kNZOmHE1LFAFsl7VoxwVbDvAeebPWb0cGTf2LaZuAf4E2on6+VIW8k1DH3/LqFTtlCGnvF8SAJQR
4WCuwZTeI8tKeQni+ekGORn4PExrbGV70wpn9ATtxOE72kJrz/7ZEOsA6BlGpdNlnA/bcsSqOocF
iBWv3YNACxwOfTu5MqxK6SPXGCkzzaCHhZFfaqpoUBxZ0uKqaO0rRXU+hEehtKF8nmcqMaYR5Jck
xI348vd4swgEuL9k/kAEVQQmegAmpXEp9BonAlgjLo+sZnEd9JWPPCfBJDdm9qAV781il1g+v3f3
CW7bnMlVPDDcmnA/iXWPzDEAaVnVhE7Svf5NsK9tTdhPulIOOyXzLtYBYRoZOLL/DoFPJdh79S7b
RzavAedynFpi2EbN0r1MT4v3AFld1lSI8PAuz50vhWlrZogLsWkZdkEUIkgRl0lWcW8OQ+Mm1cNW
8PjXUPFOb5Tf1e8XiRqG5fZSfCiP4JdLMLPbTMZa5qLr0u79UnOvB+ditDAO2a+KSvo1V7KIHn+z
rHy7K6uTV76S+Xd/PPjnGVfdXTu4w0dr4IhYp1AeNFZFB9pXb7DHnZ5w6DNtI+FE0K5IAVztjnwd
mdKY5/V8FDn7k9upZX1QyYOFx3iWi5tWYfWGIx1ijHQiYiGs90C4ECk01UoCKzBrnaIUxaE5oUAd
KLCWFVkR5SgAUwuGl+BCbq/13hn7auKWnuaB+aRxRcJAHi/QEykt8B7cHp8Q9pwXrIT1jOkC1vvc
6zKPblb41pmfnQPF5eIFKY7Q1IN9hramOBLD84eRjT0gf6DbVt9PAC3SxEeY71zUazWqwfWA8zM+
N/cNzXepUzbzp00+SQwmAuG2YxQKoTlT1E0Zsl7tl8KVNAd2x/jnKiymzZkmUG7o8E07K+zBrxkh
t8FxYXHaalgmHDkbIgI9DDnLBKlqOWX1vNgWQAooLNP3nBoDuaOSYA6CgTI64ydbKIxcC+1PFe11
RsIP+0MoMvFFgQItc+tQrybSCcg8+fqTYPXZGuUshPkzYHvJVxIm/6QKLuGQmJiTwd0QJUyHt7sR
rEGYggnednWs0oI7HZaoqB56pek/sn/7/g8WOa1boTnFKVS1pOYaadjH6/WrgM/YNL5O48J6ZOma
hJamdlHsKKrEVezBCtPT7eTUkzg8F43NBYkfjpy/ieatWFk9isa2tQI+TYLABS1dP4u9yuo9MYrd
C9ap4bJ2hBnuC3U0JYsV7jJV4vXgieWzjEvFUXD6/FbpR+jvfK2NG3prqNH/JYYcOLJcK5rmfxi2
bMglsYfwlGI9eQO3gLAhcd7UMIr8DvBEY/US0o95uAKxp/u9faXvN9FRtWyBccjC2PlZMlgkNuum
6yjAey5biHw0vZPefSUVvK2HC3BbA1WkPVUdcNwdt9N73l6nPbw6WnJkLQjpEj3PyZ6GRBtZ+/t4
cSfOkXp1LJ6AzzotsuD+H04eg++uL0nhE9GYatF7hxDtMdRrzzR73ui949hh4LnIQ1oEX1TWz8qI
Daw6ruJmKySpTttwf7Hw7ZlkO2M2pMFvGYKH0yXGlwYxdMR0eYJGptpNO51XV1Nb/eBEJnQ+2kGv
7oP7xxuYTVyIGdiXOh+Ib1x0beBgBsE7nqV/6uPlw2TDdo0o1ZJEsIL0zSOJR4FdT1iOrIs/jnsE
L9xujgS24zimLiOe5m+y59uiU2/7uj56irjh3utAnjubJB72HGGn8rEvk229bqrallwrNvLXgJke
Gwl89LBvDxi51frwdQaQzUBkQdr7nrPx1O8Br8Bs+oRXGyYfXWLksyDEzzCfUfZq1jjfKtsb2UYy
vzCupqn3vgubfw21FkCJGcs8bykDjKaLkRjaeVZ3LuXE48Q41gJNHyLcZiCIclWTcDxVncFdj5g8
Jp4hkNTUX30D+uZFLCh/FThC8snEK45tcgEyfAMbp5pb6y+Sb9eeEF00V2vn3LpcN4hbhBNLwgcO
ihjVaFawG+cdQ1LutfgibLAr4Coh6uqduc+J0fsbweB9kLW3VHFvsbCN4QWAfKbJzLGo9MRp1+kx
8Y6aYss78xgDvFm0Mi9Sn2Ek+Rl3DbVUnQy4QNV53SoDQS3fe4z7dT3lkfu0JmhateO98AoJkyt4
Y/pJxvc5WnjFoeKhLtIQReRZNGosgB2TRNIr2/p28YAzB859H9sq9O29LrqFvZXeIJVsbLJfFdjq
e/+CmFd+6bzdVfTVSLrC6EJwD0/MZxMU5/0AwFQHSkw7kP6JmKKmfQd5NdSmjIvMIbS7orijrkdk
AMaaRnP1gksgpbhXtHyqOmmBjLE1BSCZRPIS2eD3De1w2vOlwVg5R0Ry/i7G4jJovn9kXnjzberz
C6pYSWnelmCFx2oNQP7e5eH2ZDAvCDGc4XQs2z4nzNPtIQgPj7wRRXTqeWUeM57R6C+PrNZ1ko+f
7A3R2g3tyKzPktwv6d/0iY8LyobGRdfFvagbBn6Q5r87T9jMoRLP7cOuuVSSfTBFHIFZbxjJHiLG
Q1DhzcA3OAShH4zY9qwDsABApuFGLllPPQ/PmwY/xkKaIOgpN/gA8kZb4dmvaIUF8ODTr16ylrDW
Vjr5EUa3moRNO/9ABbB4w3ZWuCD7CY8RbIzXQx0y4oE9yirwV5oTHj+vjMUwvA+x9Lu1SRsjx2x0
VPtA78NAy2/6fmP6Vgn14DUt0+PYHonrGbgXJG9ADW1jgBE0tQ4Jl/uLAQFrPXJMan2eLaFFkxS7
ZHc7zsUeRovzy9GwK8tFePb3NkSyMEVgcH7xQDUqI5FYulx3ESfM9q8tqbV1Qut2+5vTuksMUrjH
JM8kvEoU8xFet31EoE2yLuFjYvfLdFKry7QTMBZdUyA5bSuTYulFPThc5ggUP1hztnt2msJlE+g2
0RDw8k7wsC9vb5Gcm5diefoPvyUTf6bB+ZFxTUhbruWEKBeUwxizGALoas4tQm/FnL2uqXzJAMgq
hkyOXFkP9FM0HXLkXhZ1REaGnUe5TysOuJw6JV8OW5uplLsNBzGbAbdyZOd2c0NhpOBNR9im75ez
Et4ciYiMx8qaE37MYkvgn8oDkCn4LMCfUkO3Mp3jHDJDyP8CN1vOe1fVCxC96DWwBbmiHnTQ1IBw
kfP7sEQKgpwtBXengyoZtHw4h9awF2AUGYeS2dl4jiyT7lHcgxf7Hn/pda5M6n4PDsuw9ZjYlFER
FNBsWukbxNfl80EXUNtD7EkForWCqfnE/hsN2EGiZfY91y9YKGDFnEQnfq90rhYXNxsnO2UjtRYo
hZ1izi7nN0dTRUVkLteyL5D06JvXyxTzSTpulH/GGwZhtMaa+ndAZxB9wAqPVxu8KVwy6w6PsZNj
GNCkU5irSS13Ac0d4mMnM1mdyHU1/m/UgTzyWgKaDW8lc9L70IyeSZdxkmrSo2eOpYGFbjXyywvW
qwipkQ4jGFWE9EO0fjX6S+uzq8xbpMvc4Xeocv8ZGCFPjy0bpbZ0ZQ1kYVJqFE9EgVSa1mTQFgNS
45f4+A6IHkR9FeEet0ENXAcEnokJeYS6MKx98zmFM0QKyA4uQAoMc6IDIyKNO+YKzocpgAV/Wv1R
50AGe7+K7GfkgsZ5DTLbzZL41/Moi6Gx868vCDKXQlnjpoamkIiA2+9/x0YnprqY10o6XrWRI/5t
pjyst/mT8T2yA6junW/KWYpBO93RFENJpG4zhidK6NYK1YSxv8U13XJKWIuvjWZN00aLLJ4vgBy/
v4gSJbrbJY6Be5ymRw2W+ArBtvOUGQniHG483/dnglHqWLZ2vMqG6vCMg3a8UgMYmhX/YN8cDQWo
tgnOsgpO8LIIJrBLP/Cye9Lmi/t3+qzB3mWpdc2NJJtrx88jBEMfJ0cvMqOmO7tYp7F7YktFISZN
Yla3UoGz2atP9Td3XgZ9duEulcQBiGxTJQvuV3D7ePo8qpmAI03s40uq9bjgAp6Cg2raSIOVVxA/
EzzRjaIGPbxtFmKbKpwMW3FcWprHrPaarq+IGqDW49vwIASlN6wHUfTBGdxr10q1JiRh2G7XcCzv
1pb4XAxX7UMrjeYyEBnkinb0VQ7RKdM4FuiERhGWs2XkbjVlyC+zkB5j2sVzxebBc20+r7iH9T+2
KfP1CHOWaahlif68oT5TE/DZTgoSWqTUPaGND4Q33lTXahJio5Cst0xjolE9TRQYtSLHUriXebKg
aE5HgeHXFDA497j5IPqV//AUs8eJIYYD8/uGDHhLZ6ZUPG6i3wk4xtF7SvDIH8mM3MfS8uaoRu8K
xNqrr5SRsA5fmnpJwkcFU4/SkTTj3XCBH96zq8CLF8d4WZfQAZivvpBLOJLeOWUwqUCw+fcAf3j1
+fx90CwPU2ZEL/n5DZDWqbUvL7eNw+C/Sb11agLYysqQ7IsyRXEXcH9jwApzAwB5jL/K/l+bg8Tn
KNbVxs21NP/Uzd2xvBCHrNUkKUg/vNidwJpmHSemGmmxp3FhMQTYX1cBlYYmdlyH+zxigdooi1rH
PqT8WvgTq1hMnj9mLUsZ0qFANV+GuDN3eBJKuTb1xBU9HmTTpElnj6zniJAS/x4UAkXtXlWwBRqe
mZmv+/dB61bVJfIISKJPWen1cO4OandJ8TD4l5X91o7Flp9tpODe7l/DdVY24jhsGFbIrg3/oxS8
sBuhJy7Vw7izAFbii4SbTkEnVKPuKTn8QJu2H+M2wEwJKUr9l8MCyX3x1jFBZjKbU1lJNUjlme8m
IniaVBSsWkJvaq8+NiPS2h3knO6UHbnUbYp4/iL4/hCQ4sIxCvmsIOMf1IbwFfIFaRzd59fKqAtD
feVughwEDhA8+Gzlf6ZKyaduRPdeA1GN/LLyI27Wh0HEqp8tCl4mgVj6fCK5JTJDdiaNGSAI7qAK
xG5r3/Ue/LFjq8MhdD0kWipbMmJ3Tgxlu/DtsqsM9PfLRqLydmBz4kYykne8FPDa3B3eXqLbjIid
0vH5PWdRz4vVIBzFfPm9GIwgrABU+10hju2TLVkU6tP2vKlIBQQsVkKIgkojf/mnDOaCF9v8Pine
WS8GfWL/T0JGAEDKFLUhQoMCYeeNGYE7zZ3OPan1+KD1ZVP74YpEUs8q6pFC5EMQhXC2wsWYxsu6
gLAKrChgvd9MAp9Q7dSr2rKZat5283D4XUN/ki+Csr1m3nSyVMpw4TttA2bGi11OSxJ6sJt/ApWO
AkNJoCIG84/WRLhnAjHP3Q+t7g5ClmXu9b46XJ7Oct2JrL43bY3Qf/+ZdcND+OvqAIUAu0KaUkjf
05ST0r+nUwgd59gsN3xl2fysdYcrMtE1T3QhRihGTZcHHF2oBX47flX9EOplMzeyNKbIsAmNkmuz
85eIfrXtkJBK5SM/sRMyS7fZyVZwjkQ21zPYOjawlmnvaPKXF2cWKdAVy9kEfWtizgsJuCrPQO35
HWJsRtMtWv9va3PI4mfP06Zd5izRmjad+S12WDT6caIaYUiTSjcxV0nbEfsnjOt0Uv+MFTGR880N
RYjDX2pw3BwwHvxkHWJyd+FcdxrAB1IFLLdZOjuXbet+1bC8CNl7JYcqk02FHtRNnHmVY61wwWUS
rs97TKaQ59fNVZSDaEBliKaKpPhVIs4N9LJzGusDH3OleHlkngUSpEaY279cl5wJkKp8oPuKoOXs
buhlbzz1SlZYZINirDJxG8o3jWFWMpBnPehG6/LTCYRSEHIaFNimyNOoQbWR42snRjKl1XiZ99nO
dxtTKmS/v31n5gzvpcVU1oHoEVEIHGCfD7RHLFdAd4jtmj67tsszgSdfl4czi3Zc+ZhhehvNjqC4
TscnVF3vRmw7dzmGGpSrscI/o+09Gj+m4of48Fxi8OdyPKTt8oxQJNuBg0s0uZuN2uV06CvBiUZy
fQUnvpPzELfz9MLOOpHpm+9Yi6OEzDXjRsHoU7isJh5EtjGwr1F1FKJ0LczGl6h00j31qN5KnJ/8
jc5kE9IPe5DokubMdi/fNrXRmxwh5G/zu8f+DyEPdAQGSOuLJ1mOFtDEZSY3kFXgJbmSiw6X+IjA
GEy/aT90WBrAqyxU7m+Ugx901xP2yMMRZ/tl6tXGm9htbhmWT3j6UA06zVFc1CBKNqJ7RVHiKipH
Xnkw9D5+29c9m/byVa+g72iDku6+2MXVsihh6RtXpOByC13AZNpFL9L7ToUP33OiINp3ZO4Q13r9
IKhondjOlGbM8NQ5RHUUWNoAXg0EhQ9GbPfJ0YeVJK2+8jDgmBBJvc7bv9vr5STcbcsksnOH/dfu
ft31ZSR1SC1MPlIpaMBwYsy6e1uVhgk7mvPAnOwQT5Ec2WSrGo3Njxywe4fGXhWwOY5grfgaHHcW
W6/FEq2Ik5wsCT5YXTM2JPRQ5BCfqmrrvDtDlOPk1AcPHGGuCcWOd6QSuiHqFYCCb0tge5U8bD1D
vLBfy8AlwiV4tcOszWWu/j4TG/yHFvjVT1k2w2MUx46hOuH1pwjSomRlGUS7tZ5mFuIdvtb8I814
ZNBwGqGQ6u+Sy8yTUAHDIMwf4Y3HX0LjdVTh2TuKcL4NkGLbmM14zvFy+PozF6F0FHB8lcvPcrB1
Y9QAwPCL8cqJc46FdRHj5Rs0C7Zthi/3y0qGshBVjuSavvQipIUfJEX0UseuKypg0KtPoBP/9NDA
wGcp0yStyIuqGhZacpOnQL0XpkJ0XyatorcooI605Ze1S2x7cL/krAAdA7DOErO9zbz275MD0ljk
aE0q+oSXAGODyAQqTaTZLBanOK7yBHNW/xYyEEl1xbf8zzNFJkpnnjE0DjM2VvhujIfWjSPTxpLK
663SeY3MQkw19fyndf7kVXtcYAHq65bWQRMXKeXa0pRhXVJ18DL/h2B+q1UKPZvOi4EhEs88o3G4
CdXTrrnBTR/JDhkBlxZPjSdsk8fdLHkFyrX819hdmXvsWA07BbNdE/tGsxoTgqgK3mpk36E3Ffzp
nGnaOF2Rr5a/aD1W6c66GXydLnX7pz9Wx80zn9NPuA55+GlNWZo8wPuQwFpYfQykfH9TT/GKSuwE
wQBAWgrcQ1VPE9AdET9b6v/IJkFEktZt8QylSFE8Vc6MM1xl1jrW8c8w7d1Q3AIoZcoj0LfJo2ms
hxDY25LZTNiKHlownnoBwiz3W3vqmCC+S10zhtvIBAtujol+aJ/oliVlx9uV395L1RgpZuesuXww
zN4Ll+5DCjIX1fXDir1/lVAquRgM5yI65xlvo+XVwWoojWUIzXXvd3zuTvajN74xL65Y0BQqmPOt
Z94TeLI2P2RRJhmNLVGPlf+8lGKzDbitPoOhr789ZYGvGgEFA4Nwb9sOoZBsv46dgLd/u94hJAUO
DJbZM2xOW7FyxkviCWjBVr0cO0Chqt8bW1b28ke70Z3GeFhi0lVfji8xSsKvW1q/GgWrEEjHySsa
xbPCEChbmCxuz7TSDiq8LvZwqo0XUdFP4erk5SRygvtm8D2MECeMQJkUxMHCYHTAzhEsMBvveMC9
PSVZHrlCXlPHMrFUGm+AkVQMaxsVrKVf5ePUnSfGdKNPP/MeS9jh4f/R+fLcXAZP82/vyfuaHirA
ow4Gvq1gTx4yhk/8IPyPgg9yN5z6P3NHoma0FhxJPNti77d3DHkYg4HQqHwnF+kwnVyqDWv1Y9KO
mSldsBpDbUSBZ8T+CsfjiTMya0V/er15HmYUYGXrkvZg3nzRUU0JfwuYfMkDf1u17d5YCO6/wZNa
F0sZ1d6dCt2LwVTi8pLLpr9xMsErwMp9/IzU1Kmw1NlDM218Vf9Ed1XK3LgJ/hS5J5dmfe91/Wq2
FvdPwvFAAMgNqm14FE9ZEH2dqXu7qpfa9dEATNHPQ+U5RcLG+a53fr1k6aH1vxIQfpiTl9IQm5hn
zW/tYtBxMvy48GeTnjYJ2Hvp3Wi4l1NTx1zkGBNfJgXMKdYhE+ar4mqQnrrylBTQzIjCoC5rhXIX
8src7lrUkB8WvH+7qrs9wTm2k8GynCiG2Qra+CC5f4jQ78PzKuG7AOoDngY+4cqeA0aCi8RNoWWF
bpODT1qQNiZxS7eS509u+2Mre10qP8znfggAvtJmFLgBn0vnhom+qyDPLt/ISozQSrhhgMkjB7T2
2ShyXvQtPB3GZqW+DHqdRxmAx/BBoI4VXl4TK6TK1vlGHZ/dn38Y6Jg6Vx4vbZCvyF+3O3NPhG4D
EUpry2/Uj04cSq4th76s+TB5dC9wIavTeQHcJgYFhooZPiVQIBJiCb8nRxsPbIPjTQ2+51d/cOFP
N1+VMhNSvEQ4JXxOzGIVKrR5LccR4RnNGmUsb/wOSImzmfY7e2T815gn/s0yJCZOsPRTh1Dwz+KJ
gtxYiBKSHZVangG7WrgzoHsDEukiByqSF3e/Exap0ZdfIguytkJ5VusFUWAfip5zFIDOb23yB5Sg
EO3xwb5nouN3k00LYz7KRtcXA5MFXrQ53rHoNCwnJT4/5X7zUzJFihRnkX4RpcLRNzFRC6KMVp5z
vrJUpwV0PwSfuAtt8Mq141Y3X3ufFLLnrqmi3u1LBWMazv5bvZyc0blAI0ZxURq1mgjitwDIlyrb
Fjho3FGHWPysL9QBv366LSAHTnpZQt/HeJbQYyDn2ztROhq6A0/i6sYOcIPFSEXa+MblD7LoQNAf
qPLkDw6C2YXcMuH1JXe4DDSQ8mocgFxHr5QchH7eYBDrGXHZKLLWeathnhtSMRirea6k5lT1QfWP
o7lSuonLupSeu+5q5RwIssTxIzfdOCIlrZkrSqomyt3lyjPrUEDfUqW65Po52Je1RWwakKgfg+BF
8HwcVUdyfKpCeJuLEldz0ot1JEJCyqdrse8RlOkYtXsd3aI+CSJVQU+DhOz0qem5foO7XhwYidSO
vVQZS/ufsVmVJuZrP5JsDEyuSiDXB0ruVSTyvRIa5QS+1ZtP+8U+Lk6LQ4Lz5oBs2lhMSQaZ6K30
9jSac+Xp8Jm/hz36JMKcbzh+1xuwPerz8ftkROor6RbWJVZkf6t2adurlDXfU+mD7U6rQ0svXnEg
z4Yso6+UpHJ6/lzse9Jj5thxiXn9nPHhU5LdbRboBuVxlSkrYfLs5A+N5oTg3UyCOaICpCL2Yoze
RAUuDucU7P8WY8j03rlq0hdMrY1ADUEcEN1hv2br9rPOoK0meAgrMWMQVU0xGATlIo7/LIOIJn5w
U29VeRRZUUtdFYkqJKXOmqTnl9k1P/LhZ1N4VR+qZdj8trDbCy4bdJn3uQ8WvYEAfsRlVM0dVMTb
cXelChY4apnq48navxbmPVOX3+0v0KS+K+dqWyrY2BgdUPXEYFzpkpGEtAGAc3yCvZR1INV9RxXF
ohcVvyqGnJm2ttkd/d+eTB4LBFkCmmKTqsWfOZdPQwnfsTpHAULt6GG2DParNgEW07yQR+iZBLgW
ukqh1o5ruOLkCRCy1BXkyApc27Xs2aG3d0tlnqM1OI9Jl+jY6eCSu46E74+oNu8LuyZLYhFVKYmD
m8Xd+x+ap+Z4a60lUqapKyUwJjhSMe1VjJHDrngTPfqHb+ZVT0M/4w5Sn8wBF3q7l6g6+VUEV6c6
7SkT7RwQOSCcfI7J5XdHtEwOa6gos28giKtNaHpCE5ifndIeK4CMS/LRn0bQde3kZ/nueU06M+AZ
iNnveToTx/9NGMRAnnbDaF1VW2A44CGFlfz5M5/Zuxv38WzefVcOWILmG85oPwyg63JYqXwoqDxb
++vKI1JQhSpWbnHW8bLFKElykSSyrClb7wgWS1dALNizUDzc36I/R7w/zIsbpfCRtFcCSdOP5eBp
VgT/Nd/OelngCmosWDzm2Xpn4Xgpta2FOoqAfEtIJhp5mR1avRDbNerSwGtim1SaF31RkWzPVXGC
h8+33S/zudy9s8zzKIqVQqpr/fqNKkpbCxi8aCMVyMHcrcK5nxfDmP9Deg/iTXYpQS0rRsDPsVLJ
mq7KPacinRFa6p9jfAa1PtP82SEBY/yHoxihpH181Uv5SjHAIikI2lQDUGn+e3cDIkMt4b8uzBWA
E5IrpVhBuxfcELYeIHjJgyYG2Fs7Zu35On44WtzXxdeZwYZVC/Jrb6wsYNxvP7kZ9EYLXvKrbBJW
9hv6Wh93vz0cHX5DuS70kaY7sVVRYO8v5Vb3Eg6Z+BrYn6TZaoYF0eFmWhqNbtutZOugNqySIl/z
ahCJIfLWlFh/o9QLivXZCE/kqL4yu48nLUrGLl96y6oCFo3hTzWaqhorhha99II7yc+ENxuyJ2eA
tyOjdyCSjnsfQleSepFCehQlGQKnQ4KVYk1y1AH687AQ32EBV8YuwxnzltL9bgXfTI2ghnp/NhNt
Q3FXBMVpZK2o91st3Chzjbfnk5BRmoT9sFvM42p3UOBJDfKE9hIKtfOZAAtxkfcw8tZDSNxnxCWz
i4P3nKUexl7I0sRm0Q2cRsywQOVAHADLYfKW/vkRX+37SnSOsVJvdzkJSjgecyjKDgGFDjNglUz7
1r1V691czv8wvvPkgen4y45L1pWosGYzEUk2A/6UpWX3uBwav+Hl2knGgLKmKnahT88brpydJKpG
ehDbJjLOtsV5D/o00eWYl5WWHUEhpvZVdHdq5/JZPmPMt9+TDEzZ7Sx21Xh6d1tRXJ4DkYRQRTTx
bky45dwe4+v2/J38IGAVU2HoFld60QTiKhNHIkVCa+ESswF3U0aQh0k1CyUvJMi8bwiIufC+gjca
MtfVLyFWTxKpEA2YKCbL+r/Vu0IGzRPqKvLocjG6NNLpZsEzcnnx1U79J9KTk6GzCqA+AjXdjtM/
KBxY57iZbKpgRVMyzRLXSXgn1mEKPiIg/lSt3WeFLE+H0shDQIxlxkzhNXZOYMNZjcjZjBb+L1cj
tCWC1zMl47paOwBnWTR5cDOuCts/mIhYMIiJcsbR1gCrOJyR7gBcF68u/iuHRT5cMHe3CpTolO/i
RhhMZzV5/L1rbwSP8HkoPQTmPBW7utuovTaUkwqmSbC58fg+6hfOfZ0M0XrGhFtXuUdJ/8eIwy88
txf1h5IO+zd4HzJAvMhlxQnqcbShIjeGysRw6J4mrdQZowrKustrEzg5pk89/7M8pVzcMdmSmaTf
fuJPY1ffzjY8TPaegkeO5q29XhTzw8e+3m/5tOH3fXVSJTbXFrcdkHXqd/2zZhtn+oMqA+2pPAS9
IBFbMOkw5MIZgrnF2Y6FgaZ0wK2G8yaitespg5DNEAkcjENaZ6+AmdfBZ92nzz4LFaayr2pwCmlI
4LtzMzfJz4MrkAnkLpjmkB8sIcIMHJP8biAgAr5I3f54wQvpx6DVe0GtoxckthNLVDvJYfCbEvic
IV1wUCrjWpXadV2agXFvQH4RkFikkQR4DHDsTKTn5PhZGcZiwz79wX4be1QFtUV/4La2cKHPxuN0
BZPt/vjCUACK0HgIEqG2VUVUIDaRxLR8+WzIFTat6MC7jL2LRPyXAOqW4kT/V8UigjOJ/+ZfL+Ug
m3npiW02w9fwO1M9WY9cZ8sR1c0lk42A2eYx9+fZ7MAwtlme39tWeEpp65zjeBblLX2nxfNMdr0T
daVR20yJLAetzyqp6pR5hPFbm1UdzYkxigD/bY+9OQwfE7ctygFrrzPoM2Mhy6NEdzkwHU5wd+S4
AOBndxoqdgixVGuzYcbtcEWrCFYGmiuo9Y7+nmRMJG50AyTX9o84SYMkXz6O/q5MZh7ReNTBN1D0
EnRiYv/mh60/cX9Qwlv7txTAB3yk4kaoJ0NTN9uM7z4Lvnhnr1/bcq91S1Vwk9LjOzUdRYDLSYEi
+bB9xDBMHAApPDF0m5+NGEj3LhH/NHEscSlw5bZtu7Xv/d1O2Nw+phPkcxPLvQdNVw25VSGo/gB9
TzEuzdoDPvKNjZtvFuI3qyVEUtBnApV7t76AHK8fTQiOyi4ueTyA0Y1Eu1c1DxfD7mqF0Dc4R/WG
dlv6q6qI8ERQGBpZAOVDgbJlXunOAOwZ6UrCiWf2/krUkW+BePrSBl2zn6n50l/pGV8iGPlkxGIE
LwX7WJrLxbYwxEqQxCMdUefVcGWkqIIZ+KMAkf6Qn4Op4yP2jiP39zZTRbs2zRKzVkceqK086Rbl
UYvn54gmVKu2RUMnmfGfaM3nhHJBFgvDqv7eGPljq8527ud6hFCgXQfKy0h9fy1qy7dVqea4fZ8d
dz4XNqjswCof94duApxwdAMtfatxBBvHEGiK3FLv+/OE1OkFxiXl6sEdqtOGmLPBNyvzaqaFp2El
vpsBnWSMGMnwxGZDqfbd1f+5gB+34NGiG8EfN4GAVv7ncxh+3xc7hg5zbHhXj0xO37s4F+NFTLnn
1lRH5AyYBbbjb+sxdGVIDnmKoYPFvp551WqHkR2n/EDHfeXWm63RSe3YYroAebOWChoBk900wrG8
zRjt2W7StGZKhSllwR4cpNv4LeQn8/xTMZJMyjgrgxyMnmQ8hbxNQKwPqnaCvCj2kcCVd8jSyT1b
CxLRgyNHYtqdpfYDjkKjrscJmkk2QHRlFHJQwD5pmbqcsCgX6dkVu860yzrywTmm5SgmunLwKRkJ
cSKT4jwPv9++ITR6j4a6EzzDaux5EQ65eAj3PBuH9FopPpIW+HtwP9cti9J8wQKhZIjwrU5OX49b
bYK80lsyHnVEtqVpIWPAkKy1pmk8XtcaQ5//oHsML5lZrmMQgOGJkAvivQXvqgF1WuZW0iHwQaGB
izJFvYU92L/QRgYV5zs/qzPHH8YxiTIiz7/5LitRjCYfauSpsgg0WGwToLYeGb8YfiEafn2dOA8j
IDVZVV+bXaz8cK9rAoy9qT/E81MwEq0nOF5IO5R7GMBp5hsTIhje+kWAV2asuqKjN+17OIjtKrup
zy0NSSuHuXiDeduJWeUKsoIbSM2z4YelTS1qCwSW5SfZa8/ibbtcY8v7rszYZIBOXjihNBKgRUln
lzvlqx1+qfvNkJ5RDTOm0lABMeInPyT2xcNRzWWSRPZsUKqnmVA5bcZ7vKR/g+VraoQX/SfKF8Fh
xVRFPZXPp2zaWvRH8Jc9urYpCpS01Pumu85C6meXCqWViKWQ6MPQzYcu0PMKbDKRRotdbVSdjXeB
jcgXuL4qXF7x95wixKcC+1+d8Si+IYFl+gK0ARYjBwHWD5Mys7YFZzW6rGxNKo9jLB/caetZu4tR
ROg6cU/i1hnYMRHSLLfk1pUbFYLqw/ZKr3BqD2gTHZ2OU6d/cQh4KSrNqyQJb207OWJsIA4t/HVc
TADJ7xBAXB8XJzkEC69wojK7AOWJtyewx4adCsaBgrwuyKgiJOS5mokSnkPiHpxQgFLZbvCLePbc
XhjCzoroWUPUeevF3ysRuVovDE8B+3McpEdIgdWKXQq3H0VvUEwDpS9veXS8BZESJNeFJn39sIqF
aq0jx0gVKFlGeYbN5s2mbgCNcjN9fbgzuhKTQfd7U/j+VGAf957cG3BY6yck9gde2Wob/X7nboFx
zpXES08kykIfvy9Vkx4aOAnmMEbMpMHPWpRqQ89t9jCEffz8l+y7nBvE7Sytcqreq5lwUbM/BnqS
e7KjlctP6cUM2HRMZUwQLkGCA2QewLtNVTH2Xbf2zYrwCX2toX+i4n6YD5vYU/qifNYFaWMSWzhe
ce15Iz5U+zIdWWhTCrjQIgzcVHcsxY/BHvDaVNnAmoH0ax1vcM5le01BwtIkDchJocjT3trArBCG
WcH7suM5DEFBDxPYNWS3Z+BOwchqDLkn048B2eTFkM8mOPOFlreetuTF/Dadh0KhyQqVXW9tVIZM
/GdQp4rl0ZBFVd2EEYP1hDvAQB8fOJ83D1lxS/kiK1IMYxxOKxJVa4eRjvU4T2t5AUzfmum9bhKo
JpWzpOOUOUHmtVz6BtEW5lx5AEOWr4EFjqW/NrOxGYM82CM/ELhuOZo8vU3g1rVvSivquz0B2igo
+Bz+meQvvNPEGD1BBwsGCcJpN0MMIvAMWtRNF824vD+pcaQojceqHR/XNOnXk/BlL7jbk06/8WT2
lPfQSoKvuAQdwtMLHHnpFnWtjzxJqdl5JbwB1jH4gB5JEkmamQV7wLg/ostm0ywMshTcs0BmTvAH
PHqIOi0aVucm+d1bfMzymi4+ktXOImlktcoTOn5xluRza1j17uLPFNI+xXtKrKfLN1BapBNTSsAB
4QsvJTXVOifhJ9bXH0Y3AROiQCF9qshPpyeC4hdNDzzwPmzEQ5QD1txUoGKSv3hbUPHR2wLApNe2
n0Z3ew2aYLZvf3+9R0OPir3xMBtbbFFgSwwLzy2vDrqeGIYDDONVzm4GuhGQ+xZ/+i5Ku1N50S0x
gNeqeZMjZ+EZgfrLNp3C14almvc9Mf0YbAZBuQ/egQpnRCj0UNfXjEYr5gbEBtjp2tEdF/LprWnW
N3YIy8HtIEhZZv3Qu7g4Ut5XI8aYfpFGon5KrAgRK27lZvHe9OQ1/mi282hvQP7ykIwJOInWyl+K
1SkE+3E0jEs0MfMjGmGS5bvNcgR5KSuFkD/aUUkJ9w8uXJeqn07x9MZWbWU5oLZlFuQ4dAyIUx/C
V5OZkCCWcQphxs214WLSaW3+Y+xVPv2GJQrFGubMO7RCYeGd9SnS9KVNW9hZAdDz/usMdC53XUoa
vMZTcZx4Jf1WnnvINVfYIjoqnFTs1w8XoAce60f50lwFGt6rlEVQCGy7kAgEVnG200/EAztLtF7r
U2MroGE3URzpJ3hgQaLRQ3uNBam/1C+UOfM+W2zuddedCkaVLyuvSYwhdH67/fMgltumKpIKVIQQ
g+AVEml7OnIFACm+RXulywMnqCWVdPbFPKj9kkUAI9/JunRPqalCUHrL76GigIoXpdERwUpQUTBn
tI1eYog5HHIYH4LiW8TLNuawwcNYSLNSKtWMNlSnEQAbGhpFiZ3pwcxG6kbbUlRNYvKyer3CxbVf
n3eLXqKvd9l+OAbOwWk0D81iX6GrYRF6b70I1f+cylTBabJZpm8FmjTGuP5DpZhMoHbOwrUe6Btx
nmT6hxRJA13IvOGkXmKKg/xV7Jnm5Dwqk3UqTWmqggdRLrFmH0kbzob5Np67OkV/nLGnoUizeEIF
Ci+7/tWAl4ijO0mFVBe1tW3pMNw8Oix7fFRLKr1LoWs8c5mJbF7a33o+unlwPSCSkOIk3B/7B6BI
oJPrkOMSUjts4/3tXDx1qytGGiwt04xf7uHCaOWHCdxZnlZxC/VfQlrdQAjm+j/jkk4Gl8cEbqRp
Box6SEeeQJ+3QLQl4sdYL7/wcx/KpLRG8PeQMvYK8wBp3G3O1JCJGgf4VcowT3Fd9L7ReM1NhvFx
MgxX+JvYytIrlyc7BSR5yLD1VnNdD1qEqTIcu60wkxYbTi9fR6nniw+hrp8N1cfo8ZcxlbD82WuN
6QEJhekeinLKKgiqL4yt5eURad6oc8sdKrzY+et9M6CRePcPFfsYAIeX4Bhb4ufjDNPm2GpTzMo+
0aIXP+pDvkTrce/89vjlOZg5e3z8iS934FjvT9XVE5bYBKTP7I1DigjB6WnJyBAV4tndwKosujfu
sJg4HDC43OtP8/y+rpwEPa3eZzoDcnlTutG9COqwGZYuGM8r9BtkViSZsuKW1Lo4K+g/yvPhx/VI
7K22g6CMp+RXDKOTUOXdr5Inlo5IlyNYeSEatqVQnZI1ilEP35pH1+9bmRXQNl0qiBMBzPQuJWm9
O0CdsfF6DUJDSZKptFwVv+OultVdKhJpl78BlyHtx1qNjPN5sEMecamG8pHwivoG2pFAwir/OMng
dV/sQ8tK+NSA2r4QK6/a7gVhCniEzBF1stcdZJg3oQiubGcg8UXPuwnXWyrUQt6MpZUasvNBoMmL
lZBYVvTJxF7nPtUg1lmzmdXTIsOu9BV4BC9etEI14Vk+Wx8ZyyXKDqQzN8ZwleUWnxN//3r7hufR
EdVXza1wFASf4NjXuNY9tkWXORAQOndFeqNkRdpUx3XJw5c/g+tlVK9acWTmebT+pg2sqzGdSEA0
G2FgE6QgWVqWGti/P2x1ivWlnS5TCeaFPjWddUgeW+B+0EF2dZM+l9YRUG+wep0hds/7mI4QHQYx
BNucSN6rkjFA2cCwslVvchItIEsfS5/6aPFwqfBNUiJm0vV20fe8vyoswcpVSg6tKQIJ05vSWhiA
a7PZAvQRVY/cTKAOAa93vdWMRTlRmmwCEDa9oJLxVxtPNFo+EmKuZopFIFG7cplmu9tVJbQzBDDz
mvuHgF5huEoVyeeDU7tzbTaYIx5G14xOiGHpwiyoTWqvtyDVSiZTJxdxMrhea0iiAaSkGBGtnvbI
CsXwXowSplpG1g/zoHf2j5S5WYHsnCfDBGmGzB3BxG9EJSy+nR+xPi6XL89mulNakK213UNkNtWB
U4RYhiEVtrxlaMlM+RRv3vXfKrBk+Qe3pstHBJ6WEgxaPEO4jL+I3f42RgY38Xgpr8WEyaQriwK8
dNDJ+WhVd15pGmQCPnKt4T97GcW9Hhmby3HheXjxsavgnQPTLsE3tWBncECtRnlTx8Ch9voTe0z+
51x27umLGJ0ZgRMU1ZAzT1+r0xaWZBVAaenhbVT+aSfPTbubh7RURMhGwwbq/aTNMlUWK2bWVLRD
63U/+YjjsyNAZLdwJW9eptGikADr9URbVxQd969V83g8uhy7nkIx/+mbETaMYHFDHm3aeOYGjlaD
yZMQ/ySBmpepwLiLVVi0SrmJ8D05vPWnypIz0wdH9Wf/f8l0nhBKVTVRsMZujOT6Pl41p4WWCQdx
52pmcqjtjTRjCRbksKxxivBTFmwfskeu3RQ+30/8iSxWBu1cANtZqBXZw4pLqjC0RTPSIPqR4zCg
AaCazPoTE0vXsaLR03E0FDXN0GfuKPV22hwtWz43ajP5cMTav2yUh1i8860cjGnuPwwfzCmbnzj5
KUqEeieGv55imt3HDKBkokxKT6qOp6miYJcHdrYnT43CG+VovavMr5zH3IMeKAtfa+tzIJrMru6H
TBKT9AQcKj9deXQnamu+XOeyuLeWa43z1rQiZ116BdbxTOaAsZyvaCYbRtg5huyWRn4t4ySwMvlR
EPreZoyum/4CtVM8gZYMSz8gn9TwFrw9dJd7BUAA+Ai3dst7p2ij0tDawhsBESnN4dl9zpH7AGm9
gLNcBgtngEIPY0ZuK9PfF46KMfDQ0gnDGZqQeBvoOa3k9qX0yde7eFCZeWnjGvx/o2AQs6rO3zP8
yn8XLP2dug9OTvGFUpTp9ok9NqJtdM00Kv/XcawOufYsuLhyr2jhg/9bbneSezxx99PdUZnmE0tU
s0BrRKIoYjf1nqzpgYffTTb9VuwkOtd+XPeP7uQINdncdpERmWvhUPizAY90edeeC5CCPDS3j/eN
/crbfcijJdJid9m0tsXx6ARd28BcyjIM0kgUcBP53yQ/SKcSVsznw86Tno+gV6nPpvZCEp1EuCsW
Is0Ee9YMJB/LrVB7GZcep3SmbeYNo5Jyy/lndslCiwGWAnm7/+C/6t7O+rnBpbn1Tn8IHow9Qejj
SlkBuUH3JGUBXmybzl95AIfoBCcMsJhKAzXZANZwbHOUa/kuIV9sTWhu2y/i6bfPumbhkxP92qtm
DpuqZ5VlkLwfJKotnvowWjGwhNuWK7ERoME9jajlEZXLZTEPTae/FgLcSB7D7sl6s9OCGk4hiFb9
NzKS98PkGEIINJO/8OzeMIwKu2QkcBATwOnZdpOB/D8w218rvpZVA+ywzmC9eaS0aFS3fTwI39q/
uepINuGrYL8fLbnx1XXqEiqmdiBRzr5UoHp9D0gcicnjXCpNh1pBZmY2OQbiSTkm8hhZHDzrP72O
lAd+Z3yps+xgje3YdhXMks44LQMV50BGB2ZXXexGTOY9tSLVGpKDILZ4Lo2jeBaGyx6MWYc8myZB
VGui2nUFuCBs1ZEKPC6QoS0mru25XuSQOXXNCtnkXCqyiFMfTVCWDtWv4AcxNfKEfPhD1xZwm9Qy
5vdExvuR65Ge9SRcSDI+FtVLAirRU19i4Q5dlbIE97IcgTeHc1T3LLXjMx8ZwBH5qnDgZYooXuAj
UZ0ezMEuQxiRFARA6aa9mixhkF1dZ/lYC4508nebBmLP0+zKQCkLh/2gOnDmLdIbS367/UQpXOcp
grUlZPs0z7fpfjwhXZgTRpW+VF6rlsq0Z+as1A06yg7IGfMFsK6t0xeNxzh/8t+ZeE5MB/fxUw1D
WAtXCWKqOsIuQlUfVAbshpTq1f17JcIMMaQqNys60yPgJ7lRlNOg/AOtKUxaoOYlW1LkT8v5LKEe
WrZdBYDDrWVlKxUXIZrBW2FX9+aMv9ZIv1kfA+tAiFa5HlV6RguiqrV3HBh/4Q+pnXxmEWELGKJe
IyQ5b1GPnCJejAGkXJ6MqcEPwbcEIATWO1bNk6lLwkwNIbgx320Ec+QGKDouE8TVyGMq0ey6yLRW
5kKB/Us9775XuYeqPET3Q899CRwSq4PS1cyymLpC/2jjOVL6BG0d+ua6Vw90/8R8wn0VKvVkny3Z
igPHqKfBFYqEVKqAhWtp2zW4kvrV5ju2YNYIuVrH/J4As77jnY8wKMXTVhLbsFpDC2su1chhQumN
1IlU9zGSnRl15HgsiB09z+vZ6u0v5g/7QDSCzCc7UcWtH2zod3ivbASSw/ggQh3UCrDXcLB9PpVG
bWdkAosz5AeNEINTcYNdSve720/nR0BYF/YJ7JpymBJkSabcw0X1uuFo8O7MOuCZ76MKC2/pTdNw
DlHYPsgB5lc8SaWLWZhmYbBn0EwhwiAeYt7aE74mdrDe6kjYdejFPkW1s+yQthHATpfCBHrFCNwm
cesw4GPU5oZmhzXq/YzKXLjKgdibVdRB0f9iY0F2IeWLBiGLIXUuXWOmA/RzwMccMZfoJ1hL6UuU
OQrlgaCF/rhPZxz6QRjd+IfwS4kCv+RdBdNxHq7RiDh4ZUq6aTzVDxvMXQa7RKKobsrxKVuh/Lng
TEUOD8naVtF3glZi2S32ahWK2Ce+p7madukNVVhVJJkUzJvkCBaYNSk1V9ZOybaZecL5gOLwrevQ
jO+lhfykMslP7iJXFe3G6B+pSPW4ZPOrGHGbVwthfrbUXaOFHT/1ID6QQNUlTtggNpXeBkhIfCYT
2DZdksWwKlxMesL5HcSW3v6fO5oljwVFjNRgD2+tLF7PbzhfFC5ASU9ZrgfghccDypvOn5nv7iso
iY8+Y441/noW0IJzFG2mZQTAJIlx8lhs/o7V6qqKN+m3/oFNTGTdaIGyyUgkniyhs+35klQIjjzz
YauZpMZ7DCO//7C5UC2wPUqd9sj3QdYIWtpZ/SeBtUOqckdM+4Z/wMdCWwmHAB7rieiZGzuR4nq2
HRl2UAAWaRWOrVb5SM3269AbWsMUUja24FCqEadNaiHy/lKQB/tYvMGfkef48oGq00mycDGs0a1M
1/xmoCCbmAxNFseQGYtnx2qvHiWICqGeFull3D+ZC64rG3I0tTfsgdp0ak5h8rdCqaBpY1nDQ6KP
iodLAxLWK0yOKQIlQsPaLvHwT2jpUE6f/i7ZUrcNPO5Tqq02th5PPlnvbXnmSdnf3/h0KMgdaT80
IKNplfhY50J7WvSPSvmpNg9cKFnpvsASjWnj9WVJikPEfah20ikFn5MexFe4+JWv0XGSGLfDVSIo
VglhWSmCIglNuBr/50Y8IJ1dQJUQVS78veIp309qG9MOWKB8+i223ewV/j+zoQh0MozR0ATnfT4h
51vVoiplvF19EjC7QURva/4rm7Fblofo2029RyJA6zpPdDdqRqB+xiiF0EL6TYSvG1Q7UviVQkKw
P+L8DosUIyrsjtJistQ/seNsN/3m4N/sTGIqc03c7QTuKiU+oAbr/+AwClJfPdK1yIChuHwWKFCn
LFtg4W6tFVWwtDom9kJhCsKQTmoxpYahUjaG1BapsG5qWZi4JbtHaC+YnOtHC9kZnXyE+ueCRH4R
/K2XZxrqd24GOrUG12s+hHrw1OzV4O1gQMoTupFqqPeLi6Ht5eHYqK/m/fL7SXA0K9JsKjGfotco
sCRhagTpSZWC5o3p4XYvhRf9EQVwDdWcJ9ddpatS0VX4utoaHtwTPMzidMUrzSLNfSlkUqLXGCK2
oFMWG1p6OlldNeoU6AX26xHmSYif4v+hV+r4Gs3VQ0lQVonwQkHAxZg6oJPS8uLtSJAw0qPiiy36
l8zevSX8zqfe7CNSHr5ild51tmh3r6mZDpaC1vCp2oWAe4G11vUDHTDxpHwPfhhOKtEc+76xDOwi
Ax9Oqi9C3btxewZMDOozdgMrLLj4rNO+j7FSxP0kTkxlovBhjLISoSSA5tfYrNCWkuV9cYSDqR9R
uyOjGHCCn0ztmzplVV8xv+CK5IqvCqeZ4wx1SUYMQx11K892+qjbdwWgpyGItAHmYmxoOlMVu1UQ
8chJKBDEecR1cZSxqlgnKl9WjUjgjImF41z+QvtvCvuytrvm2Tjz4bqq2uOmi2om/paRSOka+yRN
5rU1S6HpPEbEhex0dyODW2/K9LqOOHtv/ZVj3ob/sukeHdDtkHr/OWHMvCpMGgqfPfuW2KuSgMrS
/suI6m4Q5R7jRWunN381pVMeKE+5ACZ0zSsTyuNWRjA7w8U0BxYQZeumP21Lr/PZBqNcvq6/ESBv
Iay5RQe/kKv9vqa+XKyqAn+t75nghf79s0bWhDohNege6/lJ8t+EZS9xmtk6IQ68iuFv9AVznoyZ
RUoLjru1naZc2HVKwxCCfGqUpPTKSMA9CO3DpDen00C3z4JPH3SfZZdLPNxOutkidRrlB7HYTOF1
m7plpPGZh8e09fLUfPqtzbwlwScUaPlmPNHpvxrrvDfyHOPNVsbiTTPv9ji7+vxABZY9WjEeWy9M
bzNBC3EkV9QIqM9PVXDsUiXVRjcZAg/Cqpsd9NeZrllqjWtfmSlTPwyXZ/ew394n3Xq0Jn9qGN7r
8EIehJ4/5KhB7GrKfIx+gPwDGwbgFjpZoDX86HecCnXbBXVRz+ADSd+O2hOI21rjcj2fWrwPWLug
O17Um10zsCLvSvJ/hvK0iPqUct5LCHR8QsvaHplzoJI6WsvBtIyuNLwJIBgu64G/ra+0ylv9luQX
M0xnFXT/y07Ui+nmRtxmJZ55L+jZJnh1S10W+GqKygCbzIfdgKyJFFXthj+1JvAgK9uM2BvVkwpG
zClMxsWtG/LMPWSeTD69XdQCWUjEiFNy1kPBOts5Usxuc9NroYXjgnk62PeHfGwMAd09Jl38gWoa
YsK5ydw8Vr5vYhEdMyYJb1xLX87hFxLt0SFkFoVYCJJIAXOaPXjGaMitE85/puY6rqbz4K1H481c
eukejG94kZk2Lr2m3HFOS3jd2WCB1gSxE2qaZr03KSXbJq98ANQlfulrrwKbQY+3Pr2CjUrtyZWy
kppI89FsbyQb682ti5qYrVD44dIwknIwYNzcZD4aUzIVJt6mHlqVtrxJf/wE9xsfpP7t9ePM3ZIM
JJit2l1G3vd9bjdDUTikxYaOeBF8mesmetY1R2SKxQBGZfeuh4HkKt06k21WV5cKx89aATt1tMT+
iKYvqyrwCW1BN2Y/K2aXs3dpVEgE2n5DPHAUOaCcksM+OeIYxnMq2MKq4lcK5JXvqazr52+0y0v9
uWjYOqUlZYiJIq3ibrQiRCyNDff6mU8hj0OxGiQglx/sb3J88fGFArKU2U8tK4m2iNDUD/JHi1f5
5skeonTz75pV94DloBQpBwGCZkAbK7c+Mnb0+hsWKTCmouV1jvMvjwxkLopH4oyU1ahr5KMfmDTD
GUmBVyHkMIjx8JFNu46q41n+nULwi/7UFV4vDitgKgOvKb2FQRq2noF3EvRHCVk1XZUIu487PUoC
w6b5hy6ZKcwJPSxQLdPPzeL5Qhv8b9m/mCm8bVnX3ZRzkPQKtU+qIti3N9KCvowFUyM+Z2bBZ1AB
ryA9bmBQbxnvQni19B2cP3IKnGgR3QByOvHlN6yMWsx9e5t4yAxFUwchHGhaLLE11moK4fBs2IO8
6LEEdXmq1XvNCfsCz56orFmukvgFHjfJaAk3A5ALAYhy8OJfRWEdllQh4EjUvRuOMKTUVuwa9IqX
UQrlC3DU1uHLjkike/Gav0DXkCQv7y8zxSlLT4GO+xMkpCJc/7IKFmaatWsfBVCVUV3Ku0XoTgvZ
NMXxf8svJKVbS6majUP2NLSTVORSdYl3D3G6s9Svs1qK97sJCHqvGdpk+VSKCkj2aymyU9XzOIeL
D0ezgQQOvoAYPgvNDyOgxBWAVa2PmEYE8TWo7AA+LBhYtUiFz9ZCKhI4NJBxrMGOB4KAnQS6VwUB
pF8YSfDObvg/qhovSAxILHRA08sWHe/3kqV51sqqfwnTnlUNg/GwmcY+z5DCw4XXOK/dQUkrPS0h
XLzWyBS+1s9VVmVRFyyPUYbP+5eXFV0EhNilf2EZc0dydNzzMNxheXHge7/04lz1G/J9tPtUtoLo
fKKkX+WIeTuX9X5Mb6h3CsUJlktSelZ8T1dk1zfS+7yU748LaCz2RSrYSIqjNLBy8NTLIMsI5g0w
c/L9ojKQE0A57VIu0PqQcaQ0T1rtqjgjuTWCvJJYAkStr2xouyyDeN+VGgCdu7QRd3XDSJoL+SLr
xFmIuer59l08d1E1NTgXhdILLsqh03CghuSwSvLzVOE2e1/OSlx47hfPuityNv2fwF71WjBvrq8W
7Th+8D2beSxnKFNxMA069dIeV1ROa1XpGrKmkfWPclSTewT1e7YbT/WeuK/gIh2uHcxtVGiEJEPq
Axzi8W91TtqpWP/9uhAxu061NtddZsjrZIYw8zl+/N7jUGg5q6gsZDlNGHvhpDulQbW1axgrb1Up
wUVyKXzR+T/Ng6h/R1P45FYLSxEDJlbecb5p+l94R+GJ3OBcR+qTD6+VkJwMZC3tdqM/mkXs7czp
eJxBFBoKzcna4OTccdoHclzPPw0NUzylOjNHx47xjNlaUUFsLjo6g90NzBW2hdDfJH1eHmakkFQc
/dyZ2XkH9D79rer46dyX9pj4i/jVgyZJS76L8/yygP9eGVKv+2j07xNMWS75pRmUa+esxe6I5pYU
u9LdcU1e6SKrVsbsEh+kJ9wtHBwCM9PguHwdwByl7k2wO10RDacCMcB5uDTOkyDeOTy/QTpT399l
KxQdQqxrYC+Jwirmgb3sIJJxXfU/s+9ifOz3WkzSYsaPPXCXvivpMXTXsYBPFEgYeER82CBnlKHe
HEYfJYEipj0CSuBS0RITPkuFsiNiye7s92fnmnAAet5oToq2su89DDY4Dnlb1s48t231k+S0rls+
wo1bQjk+MKj8JPOiO7yKAieC+CJlXhCFwkaHYJrAeXqc1i+iN9CpvPo4GRXmdyfjzepWQNwZ2y3e
p6l0Dk3CJzpnO3Somx09Kv81rjF5d3s1hEY8o/BT7KQ5fBg1s2eXj2W9on/bBNao300tYgwTU7Rk
2QHK1WxFqAYSYdctTweA7ugrNsfly3WO32yBDO9RRhBq8dZk9en0SGQJBn+Bl6TKg/HXlcNST9Hu
xt7mSWgXKc64V3peR/P+ZNuPakJnHGOEWTh8LL0k9IbbApYLGkLtncuRrPjzbcG3b0GhaZcHanBS
6VPpoXduw6SGcXQCLawsvgXwJFQkJiDVbLw+rF5WopO/pl34wC2x+SvDc2lO0VaB28Goqybowj57
jPy1fc1sPNfbtQhOvm9yvegUKIn/dvXaG0DlimNGLlWp8SVojJC6dkaf7C8bSd71duylHjm36yJ+
8DaKxAQ8LsjVM37xqohppLbT/czPUEB2ZfJRLW76XKh3XUuUnBAStmidSZDJy/nqmDWOKi4a3mTO
ZybzOcA9lRxhlCNevfpvTzA5Rf6o4lWGgKAQ+79uf1TGidN0mabveNOSpih28rcwhrv0T8SmiOzP
++Yb/2G5bLfwR0HUGYLH1LTBP43Y480jThslZBiVXvM/it0B2Cv5evB5lmHN5GaU+wV9/9h4Sj7W
4h9T8RFwwUxa5sRZ8nHUm0UOrknXxu9tnQ9feHYByOgfwR+OUz6ciiq216Pn8ggbuS06rqTVb03p
K/fHcIx+/qDU4VVTFt1CYqGfWbZb/g3mEqjrJ3FyeC1F1dTEq/i21ghAfIK+tH7Dbms7wBw9Qnix
swgzhtu2+9SqBgaMsmUtY7EslbAxCiq3SvW5pkm1HQxbGCKAcKMPFLbP6yvTxobeoiuVKeflqKAC
y0PQxsA25nmW05VyIURzGDHgM3EsQj9GR8ZltL9D7z9oIIgQqtO5IZJjoLZLgua1G4V5imgbmJr/
9qV0x4hps6g1gRBdETXsMkvMLgdfWaJdDwo51nMxbKdIVDmQtLtGzWqwSrYtmOFtKrlhBZ0kkyBk
qpegrqGrln3+SiOFqcoh1w2gJugAEEb/TnONLW1M0eIYg5UoXmJcG6/AFrV+Jj+Kw1pBbHFNUR44
+nBkKeMLDfLlryr1DeaQmf3HWuyeCHL110CQ3QqL9c+A+U4gTR9k0ENmDTYn9xQKe7vTkaVra4/F
lTZVZDXjQpU5xeuhizeFcrcW6LvvgUZpg91d/1eFvpgj9W5hzokXnfkoUZvH+9do421PLX/dMrIz
WWhU2Mdo3U9dctt4KkJxTvG81Fo+cH3J7dlFQpSQWueVIaTifFrh2DOsQKKH1qG5n/pdVKME0L8P
JCyRpfUbW5AUCNZLzEKaZgNp6utdgMSO0y8zAaqw/TKKCkMyJvbKOUWGrCfuCfn97JTw2hwmjd+G
Ls6mgYVBWWmpC7XRw77nO4WCfQAocVS/cOC2UwiGJwCE1AZ8Hjt+pteXzNEIPPAEaOOixq1Tq5Ug
j7KMN+/rpZDyw/nckhpZ9CA9ffFCzkmw2NbfLI8ZemzObdu9T4l4Qc95KIARikf4cqbOcehf6++f
Q8l/8VEa9V5onUTtjSPX8nm3nyl7JP3s/EA4Jq0p9w5z9uN11IK9yiQY1u3V75ojAi62ZR+tmNm6
cBTmav/diepx91Ygg5RgSRUU0PaV+h0xf9wXboTRBP0pWn/RdADbkbJMX4TKaJd3wLJxJ4lLRFpr
lLRmjz+nPJ4TJzlhaypPY94hoyw+c6fGVY37gJt/Skns3NfjBCYjsM6j2IsDijk4s8vXsrRSWKl7
+8IBUnM/7hx87QOSrSh/VsAOEPQ5ovoGt8HLuYW/zIWGdxv5D3ocxTpSkN6Oc0JcqaOUAbLSdqTY
0z+tsiFUHDuL3L72w0RHu78pmTsknkxS+5PWsZ+9rgunHbMDckCgS4BEAt/DyFvlgAaLu4fawAkD
Va1rIa5pX7fCEJxsrInjZE2G6lAlccbUy8Zn4im1pfJjVH8wTmYvaY1IfCbbwemraBRzVsgZ/BAa
8elJNAX+oqBfUMDcJBkY53BqBNKC1savWSfLN7WgtyiG/Phbgd0/r54WwiFZhPMwyFwhSrvkH4pn
45wWgZJKWH9/elVCSGxg4Il/1Gbz7LVUFWBDcRPyfDUFTbS0IET2oU7METwPGml7aoJLBLn5kAOA
OGCQe8yWtqTPmmXbIVTbZNyneiF1mwRrXAJ9ph36KuUHmM7kLJ75/ukV7L3r6NiGKUhebhyEAHmS
5778euf1mmHq/c6xiPPaGF+QugphNAc4VeLDo4p8jfqRcQBDNpWUVjuvmoPaX77RHRogdycHQk01
8riZNx50jIGdZ6WKlPcLtOoxW9k8++GIYD5fLC2QGeZ4oqY0Z+DWgooegIawtJLpXrRd0z+B3XC/
m5AVqjibu0/Gvz/c0y5WTDcxlQjwvEml4D7I0D/5ggfxH6WmlHlmm0z825bxbQyBRwk9bBfGKW62
c2DW+O0YcSI1JmBw6Z298oS2NmD3Fy7BANEXoR0gBaJ/hOgS/jKNGELl0++ORNfr1AdnBhrAxVQC
+A2B9Mqur6XrcIZ5qsj14SAdftAMc3Th8fHO+vRcWZFO3n9Ok+xWuUectm0I24fPFLt/g4tzNYZT
/UknaUgGHBSz6rXeoRbluW6bStzQEKoVzUSWE7ZEIwNjw03sIKcwTj2BikTI+UXbp8Jf8NkjrI6j
wZwhJoQx6ZR7fVwFHM4E3L4apsfxfYnQ2dXvVizsy+8TuHijgPZ6rVnAxxYc8KUEiY28F6PUzdv4
meUMwLNI4nDpSs4HLxUNUU+cWGgk3k/aElwXJQKv5mGTTl5nv1y70bvwd+SMH4y5zmSRFmyhYBee
Aj8gZErzBfwNF7lruiAvqRiDYc1H+CgxOW3qDCOCoWXbqtW8l34Y/xhCli1uFEzq2kxJvitsrJzd
fQy/InR+CVTg1Jqxyty7TS+/Y7wvsU0cco/yltyuqFJpFrwYiqgUjUHkX5PpEKXPC2WJfSAxOtbi
J9OgKrGjVRK6rqVJOLbW9eJvIRHsj4Uvq7HvHsk7RuU+z63HbCsHZTKqbrs6uv5XTWn2kzDCfuqy
FLPu7NNAU3xPe4apZixYYHekqsw4LWOr56UtPFPiMqU42TuZU1nFwS/ywXGoXUyYLoRIgUZHf261
HA/JLxGvEDmCN1tU1kg8J3KFb/KRUW/lDL7cYjx3cd8LTMCB9XY8dnFODXxLhTuX+oUgkVpdk0YE
m6uR23KMhAvvR4PWTCTE3rBLYTkiTNPJzB5EOhYpaNcJ7xKnuwwyJFZVlVgK8Gdc+LSZ2yHqoaNQ
VNkGFzH25n1zmvbRuN5pXzk4dyxEXwC8XMH+G5uhkS8lTodpwpHVExgKfKmiYKmn6fy+DMHmt4c6
L2BvV2sVHeJDzC35bJX4z8++VO1zvIrlyNJP/V/vJ7QjeE5jPOFi6EJhmc+G7wwRZS9/ImiYRP1U
Y/dsmOM9tyjFwWCEuU2o0HIEzEgp4eqw2QkgY+O8ZSZ9S/cbnCOa+uooV/MLeywR/JqSXIAe2t0f
0yP8iulNjLclukFhrBi50j4/wwbcepHDBTuKucJOPCUGXvqPAzSPgf7rNvwQZ0lpYIsVZswjk+/i
TjX78We4GOPbbdoX38OCFSFAxfrjWjDhsVLHnQT6koqhObYONk0Bkt+oq3mUuJmc++oxCH+rZ1N/
RtM7YJO00a99beoh/tihI/EUZHKsxLDgTe1y9hzCtMbVzPe3pIIlA4sz998ehpOUdDYOIL5TM7zg
LSSGePse59xQB6xwmAnYHDQVeS/CGSLKaWJpU1XpVt/PFKfwMIXtwpLu3F/zNUzj+55HT/ajWjBh
QVr0Mz15wagYrYO0EguX7H1AdOlm9nQfw8CoQpUBELgaLP3JP4WMJ9Dzlu+EOUC1xb4CXy8wsyP+
tpk74a0dkpFB862Ra3HgTZvAJXilKda7H4ANCmJwpbYqhHhc5b7lWGkqu3RB7YjAKMCVe6pURKei
vCvS7LG9aEHnLIFRSVvwzbJvDIHBUKTG+70DgxFTIiN2YgXgxr5a9+jeqMmmKtSGhUmM1+lBrXg5
tryuzo4VV97BJpjVmKPPeakZeMw5GR/io08v5COe9YWOGj23MDW68hYhGunGiVZG/kJy9Uepwvxd
N8fzSIp2uCKNv8Naeob+7C1e7ijwgQZDK+zZ9xLcZuafH+bjReiwBewo2X2snbL5dZeBFTf5g2Fx
HAIJX9YL2UzYuoAIkd2q7L804Q52LS21x9nIYm/jODWDe7J0EM5bXdHRVmZ67Q68C3eEs1F976R9
Xn7avnpdo6u+DLFIf0dhQzytHxVlQ3YLvLjBTqYOPh7Tsm5WFTqFv2tBqLtINKAeQCa6mUAVzll5
xH+d3ySHGlwihBNoWQiC84tWXlnstOvLcGKEZoEfvWS72h0kO9oidM2Z9TTHZylcs0558nAEEeYO
Kvk/NYjLmHL5ljxMmlSNR4Z8M0e1wg7gOZ0CK8uK68o/mG6zV6vSwWAd1dYJir6WGIUqwc+3uQ1a
TMXWLtyrO5Di006lsEZe0l746PQpWo8zS+kHaxXmA1TJowg672ccvH534uOacOohlr1O8rtPrLsU
fMQ5SmtTvz0C5XXyQ53FYzPBq/JiSOYfs/GW4yBswYfPl9yT8PbLfNY7JTG2YExnNY+OEvPaJyq2
r0wVoMCLKsIdZFubqDyOZYySbpLlPqb01kqWRFV48cm/eaWre5UqNpx+tJY/XB4IHE/l0QSuIhda
FQlX1tPDrmFVrjoTqKXIxL38c/xSCj60z/I+OSOrvuPEtZfXWsnl5HIKb0cPOfvRseGVF4j4HWIw
9GoNvEwcEXIDoHjBAq4pKxSvLoSn7LmfuPMHb8sKDdiWslGul9fliTLv2Ax/YNWSpsb//T0QoUj7
JHKOURa2zwlqLMjFK6G6DOAHh3Yz2zEyl3HU6xz+RpeYy1k0/WLRQ+CuFpgT/ZJhX+xGcZf5D7Nn
rYCR0N8awkpwpKkpk0vAy0+4sCUgm9ov8va3MRX1RhQoJad9gp/DU7636dHay4IauoJLVCHvKIIb
64SUsKedC3GaYPKle4JxPlXMrEFvrv7qsx9q+zncKClul8nAapK1khBPDIyyMYL6FiNnaGwmIdTv
WF4BTiymbqCvYQl4GJ9TuCCKk3FxYyEUQVhilyGEDkaFeWy6npudu5bFKUJW/pD0ko07HIVOIulj
uijcVgBJY5/2v9jaseAggZXfao4mh574tDP1CEXV/4RT4drMnzSEtznr0iSCyNA0m3lrXgKJEM3k
7DhMEY7qDt9itEQqZM8JNmsU6ebc1IMK2UhBZktFZed9IEbfoINtO9ifqGUD754B3kGANe05GXWz
zT+2qW9KF835mdJablm7N2FaCaofLTaugAtYBy/T5/CklkA2SylIyBMvUG3/7KWBQZ/Oa84g/R/I
pfmZOXB8SX52lSRcm7fZSm6ZbIFH3IAclb8xWBcMrO2AiKu5zrAo+BfE+/8ZJPCLTt40VFNXwIZs
TuE2n8L1gD+O75iq86lHH2Tdq5a8SoHk6/E0ovm2p4KPS+FKvp6HJvMrffu06Sc8bGKV8ykfXZgA
e/RLXYQv7ml1ObG9ClX/GgiZqnd3tUggHnfJDiLCz46Z7MHcj2PFjhKqCihsNISXwTTiIxciqDqf
gze7yqH7XeW59f6CfOIX/moFm7i6Q1AavmOxAw6f00Niy15liGZUhvzqchFdaE46FIz+8t21UYPg
YHFaLwysFjnEI7A0ThUmoSPmcmtYbPRfjTgF9aR3Q2l8tDeVnzZgsLVpCpuACm0s4Zx4rl6k9dj6
7ZVwqylVce53PZPEF7sO+6NAt/QIV8h6UCfIfHzxOexCT4bd8NKkn/mGSSwiccMfQCegvMXMlyb8
/guGoi2p8VxTvV6+0J3cp0oProArdphxNo/bY4SaZBf6TtIk58mudRFJv1UDATykmfAXM0j8kVt9
korQG7AyUq4ZHwPVtgXEdkU8ID7zaE07Pw/L7pk21D78+G5xjeS0ODNCjOT8cVtGnXMvnZ1g8RWH
I5/Q5nb6ayixbJEiMjVNeTPV2Sbi0J0TWoxvwFFMiSBVQM7s2ixWKlB5APvUs3iTtZ/1b/hohi5y
Enji9l4AH9uN8PdlkiPAMUZyEy6RbFP7qZpyEHcgq90kRBbtF01iTxDFLMBCx2BgKZROqYaWUC10
lJ/WfOW4dEY98n/IujNX56x21Ynf+EZnYCgp18tiVdgicEZYjQ6lUE1m0mn0AvfIeEIhmJXEM9Lz
tNGkEekW6Rw3GOF/RyEBm74dFv9npQJQSJyLzGlt1f2CbLa4jp77DTLbYhmJcRnJsO6TKlKfnzXv
NiqZM2GEAlJLYo/F106GgDEuVKKJlO+R6+ptWd4a3jEALZKNtxCIs2xIp/pnNrzOiaArDwfbfINo
RGT2S72AWHp+X+qnUcfD3nuch0gUz/QeqoWSUuslIWuDyXPJdtZ4/gdjQNRw9T3B+6iPnTmP9a+K
98CCZjkzKudWUFeOLcUoQfIfXj955R4t33zBVFggP2TKMXbILAqBWzP/fdV4UE1xEGGgZTmNK+vE
UUNNHytMpbU1vJDbc291LYRYbJVkAWevSut3vbvgayTo4NaGge+XHAppz3nsfKP3CmWgCWlog6NC
kiJofo1k9u0C6uKNJMu/5VIrAg43tXAEkfVD/HpBPGlca4NLDTPyv7Q7bMQOqVhqOjZa8j3yvmvg
LDO5dL8vz043WNLyT34vZv4zwn0NkDns9VcN5x0vC1c8+ed08hxMwwOeBIi5kgLYOfJyC/ZB2VFU
swzJApvAfHmbM7DU+H5mllZXpEKxUfPfkWxD1HaTNMRgCkZzxqUPt2coRUYa0JGRNY1+KKmOHkWh
DPJ3IWgc4vrLS9Mt3bP10gKaIe8OH4N1JhGo/s+mJKq2Jl26FVklD6z8Xw6XjWnoQXi4eflugfNu
S9QWHaJaV4faAtgpgeNTcFnQEHKkU1IvgjqXE4UDx5NsjpBnI+lmo2xjrhllJRiOV+7vpN1i8vbW
YyWvLTOegeFiPjNskP/EVV6xa3DnyvRIJdaoRUVYOt3lU2VWPakq3IfZ02Ity3mq1zqgcfxlpGuT
qrX6awACR4m8cVpHDMwYM1cUpDllK+Ir/qyDIFKnVwyR3UrjTINcB3EywiYrdPJ18s1lhrTAyPvx
LM9CZS4Y1/3DoyMvfaBLDgVOR20q/fPmyVW9liGC+C+BJ3CjPRFFV2navIFRt7FPegJjJ8ijkEYr
8DqzcDx7fWpoq7MQs+m/A0lvStwRaCg4lna1TfFHLAmIbYLT63vUUT30UiTen3iAfv6/CM/A42iM
qCBeK2uPjaXkAGu1la1k7nmszZw0OGggZGzdcdfCvn5rxDAdDxNjJe6xPDxlfAAg3lGW/Q1TKNV9
KcH5MLFJ/YhBQNSjLrcxcK6hSf6wxzZxFOsEXBtVk14DRBG4cC5LfOaxqpxJBCYHD0fHcUAba6Gv
CmzM9Njv7QGItS7603at0ed5o6P/aPRhEOo/yfOLVsbtStB+cm1N68jmUdh+zyNLEY4ktXz1R9FZ
wn7fJlEuCSP1GR69FMoei1NpfZRrRl2jfTYgeagu8cWJNgYVP1lIEMXR269EQz9BfBV0VwgP4g0+
Fh29BQ8QMgN/i3aee5An4xMVA3zCTtgc8+htrIaRdVaJqchrNCZyErSkSDwkqA330Kgda67gk45u
SoNmF9jiJxGzYfjKBgTtm2ZyXJ6zLiFHYlz3CslCI3oNrKD9iR4Rqou3jNFZ2WfyXoDLtdUrobf6
3Dr2NzUHOqUWChSYAVj/CiMgrrZqWCj/L0f+mxj4f6K4qElYcf2puwJO8eKPpmGum8qrTf8RJD7X
857Bs6g78KPEc4udbtMQQEtv7+u9ZLfortdSc4JVVIG38fxQwFOg6wQMvuKukKfdC7jXlX9kTsmm
RY18sxk8UsNPqwgYFXlYYYsA+2FkDjyqJIXOkyq6E/MegUXH4hF3wfs2JR05vBQoAixHsFb9wpuD
KHNp94fVM6xqE0D5y+QZHkjbz+P9JgyazC4f/iyJmSHebHuymL8YzXDAljpY368CM8flBFw6me8k
NppawEXVFLr7A8f+igjVe0CjLxzrxhLHFaZ+q1HOduxekrVZ2cHhfdxQsu4bcYiVAwSY3YMjEFUy
AvhqHQezLVG/OEii+43pOvzNoWZkKABcSgPSbrp1DVTPhBENnzFuQVaLBJw48fzzIksVov7BdxeF
AIkpXZTq5gftvxvldJiRKKmFtg0kUw0JDqBcEPZO6DwWEQytY7i/hjVTXxABLldCqXyWW7WLiigS
xVC3T1xVPeRHk83ZX44EJl+AcrY2rvBKzPxzWelpRzYOKd5QWiX+gPtKQpPa6nMXT31DxbZfTxDz
7quAcjcguW9VufCm0ht6PBDpmeAEKRWJMRmwPG4aibU7qiDApjDQnGZnI1qZsfCH37NV0qsOe4Lz
ppa5Y/EeBesqqlX5bNZYDczpGsZZlRs0sh7pcRt2cQRcVksF91bkKNtyFcCrSqR7YXDerXka/UIg
62+aFzfiMG/4jrqmjkZxP8E53iYLSSKN+QfJy8hs1UeriRIhvtcw6Zbv/Iyw97h2UobHMueBFFQM
lRNafnkaeUd7BGd6wbq1Syvf3MtXvDvoAqP2snneLnfnS5Hc5eroeyK+/+i+bP58tLVB+QcmN1+y
OOyTe4fmFEqFtCWyHOTlsDG4ThebhSqPXq4u1I6aQjIGakZGKD12j1QOEdrPd6vNUb9mNfsBoxEJ
IHedC0iq6Sg4B3o7N/LsxvAyYBsrAiPDNQ5AKNI1iLw6P+OoGYvK0PwyB40uWbpDRvS6y2LBtv4K
+ehL9nvA+BBJ8tXUa3hIsQ2D8dvybqbLy92fDEcJr7ZLS+wC1HifkluBP+Pl1Ji0KkDbnYENN3RJ
vQ6Y6rZxnld0tDHaa/LokoFPNX5g64MDaAHLu8hUfDQxl95Ke7OoOfDyCFzfwuBC8fsaXhwi5R2n
eC/l0XvjFF3B7qS0r0cv5K34eOqeFiOsCd1+GFLYNl+YR/XEdEJLQSUAFsPXT/ebapsPD8INASka
9/yr+lEfiN7POIhj4KkCv7YSC4NEOw3AMpxWKBVeE7R7M3oUJUO84ulP7qUveDbem5Z/0VDuKmHb
R9/Ok60epNcUJCUCgA1TMe/GJhiC8cJp+p+hXUni/1vcyLAW0jvrbECuiqi+D6ueqGOi+PLqFlgw
92r0doNbDV7PS+CHaHpQnwjZBzoxO/WwtqUAT+YY0qZtRSgYmA3zRrSzv/imLeR5ic4NNNEdAmCr
Gaq8zf/1XfI0rqtoAI/VKzKygCa2cOK6VUwcRNSiXxGa/IAv6aEXBTH+FFtQFZ8lbaluqCXgCeVV
wVIaBBVlBT3aI+pUmDezl4Ymi8y8jtkpkzQkv1z6bgkoOeRcn6fekokUKpLxjvQRsQ4TJZgKuk/d
dHq6cOJ58Q+N3WHjOxSNnyqJZrmCMaI69NXItpf1bSPyFn6cqg+kLSwWiiQt4tmqNgsOSpE8bj3L
WnlKKZVcj1616j+nLHMBdTZctkaAQEIrY2vLRmWOO9EJYww0yX8lTANeKAW0jCSZn5PQYG8S+UZ3
ZBJ9Oj2kATMKb0cFNbnupuLp9cH5RPfLs8v5fz1cZeTf/xvD1LRN8jsqUkSpLxeDHTr14xQyvmJw
HjSYIez3F/DutTzlT6tL4znKeZ/vvgfw6oCYcwFVGaVHOIB4unDUiFcNGRvS9WscmodFGQ+xY12x
AwBCJJmPxy9ntR7bkGRN1oRKlg7w96v18Gi9YZYfQnMeM7alBRBR+sfx3noqX1KLxDRc2bSz8tdV
vN5Qql1cz4E27wxza+6sw+/hws04OGn+iQTRJxxloeTb5i0D93tjkfuJC69OCZiy/5CbtxcRR11y
nqVQimxQD9Qo1HCOTM32gTlmpc3GIsqSQp9a8x91NJ/MfGp0HDv8usrdiZ0+8ruHL7b3/cKA185I
vmXKTHFmjWKZmaVOdusha7GDwIX4tI6pj2loDx6Ok+yhFVbaEfS9LSDtfUFmdb/zfmKoJuKDhAPW
GMC8N1ROmvBuiFK8J/2RrqXiZ3Xc1+mMNvH1VjY1CZHGx3pUaHmuwTYoxf7cI8hGVbePV5p134lp
Xf2t81WgvKweSBlXhETXnAS4ce+UpqFpSbzs7290DN6na0ztke+2BDDBLdplPGJCoPZT0CSke9mr
x/8TlY3d5eZVc+eoywmORpHO8BAMcQlP5oZ4e5Jj6ij3AzvR4AttRuWwAVPfxkTIf3f0G98Fo/Pt
kq6+ioDNL6tCdpeZ1ItlsXWty3Ehfr+y1Odx8+EyFRmVFDvYDHVWeWCN9+vZX2lHoU/VxtBW5miC
7BJU5ULu1yNTO7/eP1PG0woxj4Og1wdv5lx/3vKuZnOc0VBZywt8nXtLML42LmpUCPIlrTnWQmfp
PRQRDHsn2uYMoM1hYpBYU1m7+GhH2VI1IkNBU2ckyQgCpE4MnQOnX37XhpXOj69JkNlvs+qbU2Po
ejq/PKN7b1tZ/UTW41MZZug69pmD3a8aVzoOcf2QdskscEBxKSNqiLlVXjCL9U7JvrHSFH0+1ZOr
3R766lfoLKEIOwX7lFgLa4HBKJrmclI4JBebtVb5AOQUtPGVHDDapOIYMjneel9x0IvbIGwWOSFH
BjMp4l1hDZRTHOEL0GJY2+gdvG/+nq17xC8R1bbpuxtOP+QmLbZK5EM/A2g699vdTZAxo5AjKYTP
98yhHHCC0efR9ZfOW9Hti2iuN3TIf/ZKzmjRX/IQMfEzYj3vqv85hsfHO6eujPEwQduQL3ZrEFYH
zmUKghJv/mS/pDSUgoG3NqihXLqpgyfgbv6hVxCy5OLxmn1IY7z3QjfFq8f5It5gFAgvoix4BAfW
UP2UqF/+jkr5Cko0uC+fHLMsSX2b7x7MmV4H1mDnTvDpnXEbuxbL/RLq3IW+/f2DhOFLt6Kukous
32SADZQb0SolgzBoI2b5rnK2yNqrtxpADb/TYI9bjLc3Eo7P3WHoSOqDXsW/HiJRCDrQDu0ta3sv
G6aXE91vcXv+FEXxdhDucpXw7wz0B2LlBiZwMv/Hep9cSdmZGPu1RQNzkolCEUHIzLPa9KhrwdaO
A78fgw0l5rg6uRbJzYvD9Ui5aP2qdLP0jgrBRhmo4SnFHykoyhnBNEl2Epq6s5egjA3XxHKnckjJ
Re7HFQ4+tEU5btumf6sBp2cFQef32MySheqkSr2uWbAoVs1nmJMDfiuDXUYrr6a4lp32Y3I5QRPd
UyTWNQkS2G7UknEASCfurbpAau+pZrD6awQ3PxFPBCQO/z7OgdHFWBcPLi9eCBpWXub1CJ/2YmpD
gVydGqSnr0rVQWIPA/o0mzJ8QidfoAcQdMlHrs9sg7TLptDeilaViWG11p1JafDzTeqAsJaBB8Uk
0ITFBeBKqr5PuO0o+Uwc//RQKIvM3pt5ygsrUI2LT1R3YwE7OtlWjQUO+J76lFRjNU/tiFv6lMEJ
ps3iPRpPxxSZ70qk1qi1lGyUPWIp/xInBN6n9JNdixCMjf73d/CLkLtdf8GGh+2utG6duR/Nxa/F
Akd7ZG/5BjRzFZbZrbxHUETopPSDWJT66zgg7Q/hqbDxcz4vBy1DWMP4xM0tIt1M2Kqb35o3z98f
W17CoaTrUTFN1jm1aFdm+JDL/uJLR4vUS93nbK12MqoE1vmbtkdJV/UABng5RZJ+PgG59qZfHAA5
wjSK232mwDGMncz4sXmEzo+4h7wEXuRpinoXasKemvimgK81rHFps81+lFLNbUt9x9WVKl0ilp4C
J0FegiCvO+9tf8YY75t0HXsDYVLl9f+Ee98DI3FPdg9Fkqy87CxcNoP0LpbrC+1qm0lnR1kLaRqW
nTrUhKND7tcJC5w7tPWMemA5Pr5jIInm/Y29ggYnTqW3notnUC4hE1FHnisu4eCsfyzBH9pT0V8a
oa5gtnqaotEbnOLwHHyNhMi5m4CtWJsgmcdZDCUoSIEtJYQLqwcLxnA/tP2s5JkSVJOpXDPCItHD
JtpjWU51ES9hDCTpPb1Zg0UqmbqiOTe978VIQJ5woeqAW/c6VVJeXm1tBGxClnGrakTqjBJlYw1Z
Mlt+rOi6uixh+9qikykwhE2JcHcQBB5r3gg9enyrLARTPDyYk5+yU/kXOKlbnoVWx2xdSLGoCdfl
ks1lZBB2t6xzcVj6AVnqDcIoyBfmwc4tFo06tepPrYjJ18jJn7dcwNTXRTEiD3ifmSN7+1IzdVKM
5KGv9J9/Z5cSIkjXS+LA9TrTzM2eXEeJm86tDrc6dLxqGeM99wijC6tnmAsIwuqq5eKEZEaX/KgK
qBwzhMlgmnWBdQO4ktSIbq+ROyFeB/8iw5aaduK5RQjqhXOLy/br78qfFqM2wH6cSqPnRoLfYa8l
XocXN93ddX5e93AafNIsAFPD7j8ISNFsDkHIxT/Uwyv4PHHzx3KCn7CUH8EKXOoYz6ueSKf4GVFR
ffW+5mxN4HFEBFcfJ62cQ9A5rdKxFTg/vMRZthX0LSvJ8F3159fJtNa8ahi1FfvDFgPoOvuFPReF
e+O6IhGI1oD17Db3ISfdv0nhZ2Q+uEyqpoVaCGGtgR6Uq+rz5p5P/7O16FVeUujLf0QrKV1J2yW7
1OnU8WHVncQe4MPxYUYJkgqFDYykHucGM/ASJfnoGb8iRm1V3IKPJXKM2wPiiCrIGegt8UFXjMqV
7TQn4U1f7G3gLcN6rQ5fLBC+VWIwVNZjlvQwa0y6TZsUkSSgoA+f/tyNNaV9WDfI1W4gaJm2vr/p
KDLGNINdYpG5ryZNXvbiSHc35UENsx81x9GnzcoEzXHzI5qc6DuT8pJVGuaSz1p5AuieqklLsjMW
jnca+zpwIUsWBKrFXzROu7VXVuMZw6stiol5hrNF8lFRWpJGK/TtXLjy7DWX7S7o0pHhKiM1nZB5
iHBp0W14b0mm+jqir4ol6nFopduQR4YgffQYc9ag31Ps2UZc6PKy2W8mvhmF0f2zg4p9wAF/t3/n
M4SajKh3CWajWbGCJESmyAce6/IHhr1QisJB8gMtEOJk8dt9p4KplvoXvvgNwBoP1/szoOalq1mi
Wk41ucoMu0Dkz4BWK6ZY501AbKi301AvFHCeffzutiuVoBV1q2s5Iqi/st+XsQiCAbLyLPOvslzE
fIdCb8dOuBxvSoY91zvu+9GALs+OZfTfVfC7OYiRcpITtRIUIvYlRWFL3xORPSm5LnAM4bWfoCuD
bOxa86HYaaSVJHIuebvN7uKStsAbeZR6OLyHKTtuUL/QpwxvpBRcf8R9IJkMFnUhBoBvfnDKRo5Q
cyPgzbS47qf9+32/UarQeXZACgXv7oKCF1hIIPW+UWEQtWBYmkcu8W1K1plvkkPwjCpTHwerLEMt
BZcj1jJy+itJGH4/ySPT24lxAEOzWvWHpak0yONPC7XsBjFVx0e0Ctaxw709HX680HpPIX3oF7Do
h6DbCdvjcwH6Y6aJLhilk+JGD/jCYwoMyr4/1qfH5yd67I9utYQleasJlv8ya9gxthjHY5mTkhKy
9XN/fSi7tfobPWeYsZ6jb92QP+Wi0RoayKOBPuMFLT77UEvmPk0Nfq1VO4mOf+9WRxzdNTDXAUEI
+D0YuvAuWOAgybdEf7VXvXeylqxORpuQ4+YNpqT1gZ43qQeC5V7ksSEpq7EJQepeCFTk8KBlHamb
7tl3PYEqkP1sMz8hRXPRk1TTffk+i8V3t/oSykky2B+4RIMRnTX0t78UswD+TH6lxbQClB8NxGTg
HQqJ5iqcDAD0U1/fkMcYdSyRqZlxJkjYmQqBwOYJGAxqcd/mkx3E2qKUB9W7U07czlYdCSsyJTB5
WBh7gQbAme35HJMof3VX7mh4vepV+MiO4b/XaLLjsnSG14pObe18QCfwsxoaO7LTw7If5fngber4
e4iNMsYx9Z/XwXEW0Kbaxs8ZWi1U48bsMU4anOC0PIwDtxDLqk9PhNOCeYkyUsdyShp840UslRLP
zKll9qKf32EYtpUhrTbY2ApkbqUD8cJstiM3uWdes89lWZFwrRv7Y54TPZ6ghqEdAJpCNhfdHCFu
8XVqECdM1P1Dc7dus2M3uoUjlJq04zQZ+SbTsiw8mQeFcBDXzus722Y4YfUHs15FL6xnrO50qOY3
UPZmylK42Ian9L8n8DN1GETfwTNqrTEaeu+NXq2crIsT580CWxq9ZiWWqIouOTrs+9Ldw2PFQR2E
mQ+locUaVidSszWnPCXNi2Fhemb3uDB8FfBZpKjzkRmbcFELPZVVUTa4CzpmaMJlI271Jj1mrylF
9YFdJ4DVTfk6S98VoY3wWS7v8VLNcXOAaVuFxM1mezrM6rcnHIUKSXxmrIvgzBHXFJCE8Fh1fT1z
MVl7vB5dIlbTIa7vyGz77VFanjnWrUmzaETMDjNgz4MsRYQkSc2lUVtTa666eGoAzS7vqmQotH2y
3PqQcx76TFkSmjhZiweVpRDugZ27w6C1IpIlPJ4fKXhBNp7dvhdWZ5L37WdyNMdYvKbk3PvMPQjv
Fg6kt1DM6Fx/1gi4OF/96s5HigzRqx9ZmxjR/CQLpZxtuHXouIq1UsfevaBxlmukFmQvN5atMpcQ
X5a/ixtgLB+gvvJxtxDmh6xQmA8QWR8wRj+d6CT0bCfmwUPhQXOz1WPRDk+XXVAfvAfk+KA6R1MR
kmOdmNHH15LAhpBvKMtgTnqoSytC7bIQqz3sYPtWR2QKcBQhg1YVCNQbMbuZb8LAMYnxiSFNQzFD
EncoUKMvKh1bN84tgBZkQupGABT+sndy3REtyp3OVf1e6szTN0qGk1ZV6O+vyHOI0/XQvjTGH4/f
QhKtTslE0g+b2uIHZcQTA1Y0zICjIKvA9enaQkmVHMkVh6j1SkW3lAnZjqulk84B1ZcDD4GGvwu/
9MZehUbN2CbUsLJDWN4z5OzgMAE0LLrJJK6m0/1jSB78UfQLJZuoc9QYMUac0SirAhoTmMVZecLj
lIaop11/QEYuSwwgOJ9P/qDH92YSts9RjEA/udymPWSNsltGwg+VfUvaWhK1VajT9iA7axeqZ3rk
K/JyszOXD+LFcyJNCyr2PZFD6qh5vxgm6eUsPuY5r5Z4fpNglTRDuK7mmCfRwJeA4SipvfE4SKyO
d14Dt1APEGqgwVDt3UnRQhNQLfsdX261kjwqRK2XdzcNglTLlOEAzmtOwiFq0i/UmyzRrrFF+S/D
nBQA4VF9bXfoisdB7E5Dby9SHZk4IZzYtpFJzNovxG7QInH7LSqs9qQKIc5ZN6hdgIUoc94udsLg
LYyxv+GELUCvYslisdmpyymzLZvgms15uoXZj6n6tRR5GVUymmu8ZBELTe9GSN06XpCq21OxGmlU
inRz0NLwJCoEA9iSRF2dK3C/bm6utmEMjS0NK3YhAkQicbXc7RPvvzB7fZgDSxilDqw3cwvlCxd3
iVFT9tWTagC34etY5Ogaxv6hjVhILVFZDhumW5ttgdokRXDywFCoujlK4nh1IHIXtiR7Yk4OSv2P
tuzS6U4SMlbAPtcFvFLVC/RQgXXJQWaQd9uidgOo/bAFUgcOJgRaWd7YKv+mmN+/U/t5Tb1PBhef
UsedrqFl5EA5AurZT+XmNJBQFprgSGmPhZwOr0zmyuzk+CHkGKelX3/EkDk30xj3E+LyE2a3O73j
CfOU8BtNXNMfXLw5O/cJZE7Bq+r4Ux7ZXaxwec1KrkmQbtN+gaI+qUfQ04IvRPBwlZCda0qL+4W8
Iv7G2ibBM4dYEP0wYbLRaNgDFa/jFlurb3Rlp+vG3x3BH3Qc64ha7UkOal1KDTW19AvCnBjbhW9K
PLDqDR9yDd1yImoOGUwc5PD8Qyl7SWnEtCkDg88vWnJvHK1v3mg6+xrOxRdxxw21NZZ/r8YnHGhR
swoHHhrEAihpz1DL+9wQ22lgIrQTdz/70y/KDRHfsU1K0QRMT01FMeVFhOhJ4/Psq8hRN4321/hz
0Q23Rb5PP0oXcrIpx7fVy4a1Mxd1pMluPsN7AQGnV54MukcBppUXhXDiGz8VtmBHPOHPIwXwVJmt
FzypE/a4xRRKUHS3zSvjeCCpurvyr+rEJMDp0upa3XLGp3mi4XY2Bxbm4fQYrtBoVk+elb7RX1g3
xRPo/ngCdPmpAjaduyKEeRdyjCG3cxMqgwXSIe+B/XfPnYL77KsM05h0I9m3/9jsCRlLhe5IfSgj
NHblxIWAd9+C9lba6wMitYDKxsuWaRGFUsAoz/Gm3dKpN6+lK2ZzAI+3RqJH6h98kEysXQQcbe8C
oYTbnyYkhSwW2FoygWHLOeQcAMrsb6zH3NjjF1qx3vpMsCOGil+CmktcotgXcR8nPDwQfdVEaWb+
kidXNN6whFKnYfK3MFcHyk7csmiMlmKRShT8Jt5Eur5Mx7DkRjNgjJesOvg5bcMDtzovCH8VFgyj
rpqUUH6wn386lGN1RM+LIFDOCvsT1pbnuK2Y4OCPWuLX3iODuqeQGhTo+Gkdb7DMcS2xCB4qM2l2
fOx3jt3UHFE4q7KwS6HakzOOtMXpdxOrV9SeRSVUbgYv8zDjbjH3rdKnB15e+dW4hOF4rseAdCLJ
EO5SiLYX5blMBcBzdBbigAlX0O1qaeFZYIbbRkU3e4stKsuEx+AMLQBVr2Z5xlots4GaSGEiIhD/
+SNoRN622KYCmOx1geZ/42TKaMBDmQpP+8BMa0Wl+es5KLzyCqNN4ofp9E0xZdBepqZPPu31F8Nf
JmLIq0Tff9+stGnjlnN9OcOsnLv0tCs0ceRzSDlJQuu+pLXuOMjOzXsSyanVVKgHEAcRFfv1M2HJ
PBEPTWdfWhU/rC42OjesOk8onvPCshnyg3XHOBq4WnvIBMCHkrfKHf63EICT7uXHMMdlwko4TpSY
KG6QpUTaHdx/H4IARp+LPTgFQw8Yzjb7zBwrVYTLkfYPRx6qucNhRCFiSwmfVu+WxchCeOjJjqnR
CsUJGUPxVX7lYwl87ZBiSKx8mCbi7vWImDruKbaKV0P03WNH4scYSUo3eaLg38wn3b1WE6XEAegr
GhhAOKAzkZTwZ99xGFDSynLaRYh6uant1jP1YIfjaNU2oiU0iHTgnPbpCr7Bqw9eazcIh/4vKV/u
snA5EGrb7ar+JKuuPNecRXlGvhc8FKC/qfAiWkc6b5GmvVQPYwPlSTYYDgENEWDnwOJZDa6fDQPw
+aqqPQ5lbMvFUttVjSJYwywVjfj6OFMOy1uy6MzZlykELym2afHfm9wx97+wFhaAmqlOtTFp2+Iu
bt1auZ3xiew2FEFiEzMlZDUzal0qvTkUiKbtra39LQb8UtvedRhkLTFQGe/MVAbZ+MsCthkrNDzV
c2C9raI9SCNN9OGTwKizpAlDvOYLqX6lzMkil3FdE5yYgun+dtwjUVtOd21GEWKKkXQbH4a/txYA
YSTZj0MryD971/D+MAz1Uh/wAJWDwCMayimu7ISWPU9lDYwMSenops3TCVTULAoCYUgIEiE0UJf1
1dGKfSnJ6Qlob/qUcdR29qOIxgRgJr/eMRJESR0/pe74o25a57AxJEka04J3jRbecgpfKsSMszNm
nA/l8ze+FhZzue4sO8kG4yPprIdgmVoVgFjgI3eGS6UPReXDGt65TPZiWdeN+v67Lydb+LCVd+nn
IorUq38Ef9Q4Ze5rA8Zexr3qY2pX5YuZzqCA1tIfL0RE/99TPspjIkxhiWSqxg31DqayrEDZKm4k
2ctC0KrWZAssNdt5cUQwesD9dkCIQG21NTUQSVKUGJfz7xzrc51l3BLCb3e+vw76PlbvYXYOGRHC
k2QaTSt5rgB44jyRuEbZIUbsTiuI3wkc9l442NPkH46xCx7c3+maW0p+7fp7zOl0bP8mPnVvYym0
p3wtT6PE/UqqnlKDf3JsPRVxf1Zg/xZzYjiRtyojZPcnFBYpI6OnT9aEiE9J7wNFBj/a20viYjPQ
lRtt2kUYwrvhbdXjEsfJnBClXuZrWRLPBvmqQeHNM1UldN4npoSfLPqR7TPp/3g4+UdKXxqOVJCS
AWMtmvG0hI1gO6y4tByf8wPgfngIOj4em7Unqhax2NZvhqc+BbBP+rzYRQmJtXu9HrY5vlufo2pH
4f9XT2S9HQ15pO95reRyloCnZ/P/aukUWu8MhQprYKL3WdlT+bE/nqw7o3DWZJTlD9FsYIwbG80v
/9aTcG6Kg4iOjzENoyoV6dUbEkYyrY1uoyTJxFxaXe+ohL99PIoY4zxLeJdbKhQKkU7qKLWBotJ5
R+BnWBzQL3aK3WyVNrMXY7RXMhnIGmhXO1hcoT09LaT2CL5t1GlzFE/V5GcyWqh+vw2VSCRyaact
6a7Y0t1PKaIJ73oEhuW8vJ8V0ztvtre2N8cZSU/HWITZP5cXlj+gFLda9gUxVwOdOHKR8UJQMR8h
XYu8AMVb7csrL9ETdKDGmzrgZReA8Kv7GdAc5RYzwyBjlGLLX0ksAdYhSZBhuB47nvpoJhQNqkfY
JKXzyyZ7PVw+1g9RIj9zQY7HXbzop14J4X01cZj01NSU4seLiZNyCS+QYUBbjRzvS+lqZLv+Tic9
3vNWnb7tXfBQ4Ync6N/yw09CXvqjPvcoPmFnLCnNtevVZ3Ztos58qVdp6aPhOAjzn+zd5iE406ho
6QxxwherhjFwpKp0F+OjcaiEJ2woMmLwaBGBUy0uFCqNy5AyngZuC/2YTn8ffdBV70/OED+TTtz8
qIO4EaVb6Txm3FR2c1oFIYiykl5FDOOIeXo54ObUcyq4ZFoSgAUv74VXCTrEjdywsECuNgXxQ8QL
UrIBjCHSmXhsi3OoQRp9ScmzRiYsrdTr2Z6NXf2t0epb9HLw5p1ApyqUnAv0mEEGu/DHqxsMf/+K
H2LyqfyRCqdFm8UrAiS0fMbz+uach22uYe4GnDa71C1JBymc2O2aU92j3NJGW3pUJJ2nzvhP8rn8
NrzoiKQ3TT/fZwmPmiKUo0RH53B394jpJQaENC4yeIInmPr/2h1icgw4tiFI0Qe9OEj9oYDwVxKZ
dAUPVH503WUlnF7dVdKyZnlB4SeVYq3crFwax3XrjTkLzTCwQOQFrqMnvLPX8t5gVWByX3rSjE1n
4cAWol0Rb9Df1pA/wtqQ1FQ71UQngfLPPHxmmGi+QyXrGaIyIGSK9hTq0Fyr7s+a0WVtVv2/DS2z
4dpYb1Its5G00+7lZcdG2PVgDvpFT/WhVFjfY761U8YPihc1Y9TyHU3rN+RDxLOvCQpnAKiFNeVy
tbtdFGfrKdwvEUXMd3gHbywKBLV9naY2yCqSROorxwwLxPhe8NGZvgLLmW/cug1p2LmzBa8dAUuo
yUZ117gNxxZP/FhRl3+MBCetyRO5L/qOI3QGYfx5Ak7iKoGC7RcSosGpv9FsAOamPO7RZsvCJPYp
WiR8McSglY/Au1ImiCC+0AQSQKbXtLYhF7GWmG/YPRhxRTKV9smO5JDB+v//45LmLXYDhvNE6MxT
fbjmuk/0h7lGzpePK40zlZRjoZBieK5HP8bgZSVB7W17JLyXidXhn2Pj6ljZ7uyPZB5u5BFEz663
1nhKEPXhrvzqXss2lC3k/reeoAcyafmT9+80ij5YgGugDjV/vBZ2yqJIR4UFWX9cDUvFxqq1HIRI
sYXCbcblwNeq27vbWWfZSDTPcYIn/m4mzQxBWE3eY4LUTceacXcZe7smUhYovLVg8JV05F94emCk
Z/tBxZg9T4+AxmK5lHNq1DY+HMDAKQigijoz8YWy4gykJov+byse3zjnbo9nWmTRz00yEd7ADUWF
fvGEHNaMcbHH91nlU2cbQU2pWurAL1e6Q4JKfdUjcjOjFevX1PdA+D7xCbbAP4xJ51XRaIedlT5A
swNEqD0H9tfrC9a0kiDUbAWJxREbkGO6vanRgbRwExz5qY/ROvOLpBUP+ydSzb7TteizXhy5Y7JE
NmbkIPGBIZcg2vD4TeCj8QvPlBWwCXJVbn9Icv55GH5i2eddqoGZmwMvWv4uHu3ieo4AuE3dTfz6
LV7nrJjYVxQpI6443e5h1frR2a0cDPHLE2XJZ26yC+jXgn8W1pHuAIz5J7piVUKKsOfxbWMq2+EK
Eccej/UIW23SiS8AfspqmOESNDsONdvkYrgRnMMvRaBom1b1ycuoDDJTy+EllODuph1jedA0Zoha
PU91F8kAHwE8REbjSZTtrJKTJEqooyBi4QoY3A3cJ52OP0yQZdd4BPrrw7NuqRWZyEfi1TEYktXk
VHUAxnU7MTblNCjkqODFU+CulFgyz9OITb1UQlzLftfqphmHnxtPMxiAUGmPlM6dUEUR/gqHRuoX
V31pl14R43NfpqDr/bAk/IEzmQE/uN0rP/ZoWA5SiEs8EKbYPkDxqX1FqWcVcOFJUOyn2Nd2JUlZ
/1kPkcQA18pH5a+uAl4KI4BJjuZA/raBK0KU0W/BbIaBSw/AE/TfodRxdVP9kR3wqhLg/1Tmq2VS
NyAoATwlN+cxXSD4HV9MhHWtF21yGJzI6qlmBJb22zIfoZtD0HyzBM3x4RH+2WUmOHoN7XdjoP+T
+hswVXhZ3pBR6drvXXWD0+ZJozvGtbibX4PB6c09XW622iN9lJgT1R0GW49tnS96uyZlG45tg5Be
r0AsRBzi5dMoILdqruCxVzgPgV5LNQ0hBNOxLmlJA9QjbNKL4qNuxxcGynAJpEAXbkKMVyCCqVFO
9lOOzjrdvet9y1o2P88QugihWJjFj+jdN+7rU62yfhQQAbc19Rzf2lxANqMRsWOaQDvuRm1PiLQF
04iv1QFFug4r6lUwvJOH97sjK/Qe48aGoxMMJ7Hk9nDbo1mXrovugA0Gh1ASPyON+ARE5ud+IC2Z
ttVUEM/LbFx38i/DHU1yDo6W2vNZ4B701oVyyclCzN6Kh+U6P5paVp8h9JC5ffx4Gc3n9mfTCkOy
xfkPwdIAmvlQEGOxVOciuwxbB5vyrmTPatSRBSIXt2WFnRZ1nWPD1yznv9lPgfW6zg0XWzr14Rxo
CJQr4P2yHxt1DqsTsWvK0dWDi/GxPe7W85mAp7tCDGDtkYhUkXpRtgQ94h/tVkjBq0H+2oASvzQ8
cRJ2QP15zGyR45C2ZeKCgelTOON6LNJ2Nkm839wtImcfRffaxzhGrHv0eDcf8MyZg8dxNWj95w5a
EDigQmTv1FkL1mkzjdqd+ZDH+JJpbipnIPgeqEAyUbfR15OgYY3zt6nJDCiwsuTGQAxDmfRqD2wf
3E28WAs620JcEcegiLgYGnwlMVcyN1WyQ2cEDke2AvWzwobOAdvjYYPLaf0PLxqT4aVA6ga1dTa3
qly5MWqrVlR7HbY1li+swWQ5Wv23KUVVrji+ujI6Vy2oJTygcMoqZSDjkQqW5Lkfzp7Zs9scqglS
nFHwoUf06exG562wzHIyKuFUSQD4c0ix9+nF/Gqj5Hg/WX261571qT2YoGJ+ezlo832NU2fOksVW
ehevJtL0P0HCd5nwT/Ee8ostDaNID3quwsdNMize6UbbGkBpr6e0sJcWsa9OzX9f8W7BajyWkjLl
xIkrLBvvOQWiM8AM6ZiR2h+80qlYkea4H14FEHQtXeTHmZAnk27+dHmJX1bvubGeZRkcLGzCzB9f
KDevLY8czwkE/3GRE6CMh543vzUDdQtxgPZExwkaE3FyW2roonD1Mp3+QLcqqi477ofSO54dQNbv
ZV90PqzHa4Wcof0VJ13jSpVDYvqR9P56Y/dTMiXALjQNey30RAIETWlv8aCwHt0luBo9nZTqI1YT
Wv2NoWR5CXbK4taH30e8asJ+G6u2fGUIOEigUQybbGys/TmbEhk637Nh8RmGIEncq45e8wPI2yHw
q+Bw1XHmua+TbTY6mRFT6BlYaltROp4OoJcFUwmRkDt/fNoXVjWquU/HuVJUKTl7JUmrPG4XATfW
s0zRYkOfsHjuFDEv/MwwQ4KA3tUr/KihHKLkpaG+j3SSG/wMHojxiKUmrLI9DEuYOARWLyWbPIsZ
KYYzHLydHsjH8dG8PAVnToL6uy3ZyGRWhuQho6wEWd8Zzl0QqTUU+NDELx5L+Tdrm8Wm7CzHyBxn
RUU+iH3xwenYHtmLDw5ELMxNyfDJZnbhbS3K1FVvl0BRsKNKRluF+Dyijt/A215j3Dw9wzziMGib
8vvN8SC9GhJxB+qgzsNOFWZjXTtNfZUG19bXukk5s/Pc8bCh2WCihGJ/Lww4qjqumEhk97OvxJ9J
xeLFNhiDMbJOusbnqVVFC7mcLwDw3y+TlLdcvhOuc1IBp1CBm2WEYgbb6Jqqyh1+FOi4CpUnSll/
c6xwnKMaQ780lK3UzsJpmeyaJwp0v0mqG/6OTZ2r80fiqdMEv/Hw11Q6MLIaZC6Nb/VHODaFkXom
uDu3RNpoDETvSxr7agSIlB8zjdyziRUE9N+eMr6a4rXhXQOJDOd0Xl6pezCLyLc7uQXH6YlsdWBj
sjR1rNZhYxVnSG+dtnHbZWP3vjWh81YMeTHFp8Fa9judSyYyaY6Y3ud2MZ9QbVU3QD7l5UQlvgkr
TN0qRMj0w7hdG+iEkWjd5B5UFM4BClEklvB+wwBOvguasE4Iw+/+FeITmMxSNQDWq44mTSOAr8nX
lx9vW25vMpnT3m0sTWglEzkOpMsiD4n8kCKodWZb271QxUXzgazrLTyHR6ssBe6mRRMXy7CdFsHa
xXMef1a7xrhgjQAv94VY8WTklu1XfkgbQHcYx5wUwc0iaUk5fra/ILXQnlv46RPy9fiT73lQEA4t
Ub5QcZmYVpXBcJm/G2Y69pE3UOR5zySadonj0/VNOQ4lXlHj+RXvUhZrPAeb0YXm4YkNL455pEpe
uy4zBPMAAD9jqTHCcjZjAF3TNKIFW6yA0Kj5ftDMe+EHMwK4c0M63Q9oP7JhEapHGawKRorDolE1
aaku2gmgAJEA8bAgHZt82euIoBYVuDJsFRkAfbPx29ij9Vbz5//5e1/NhjnITbtezjx+PeoV8hDt
VwPTY86GtkwRcKfKrzT5BR5vxSAQwMDk/3YWuaUmg+gCNmrlWOItZzBBsLz1IxSnkPqMz0BCG6wR
kmQNNhMwJuB5PTGnIIEHbGUax8HNF2C9gA2B4+8YcVsn6EOibd/so6t67NVAVeJl2tPRfW8eVvDc
lfkpL3+yYyv6fMQmvi8kpkaSw0tNfUz7GIAnRsFz0yOEWB4auQd0BfeO8FuJi/9hjeaIrFxa63yJ
i5Jh3LpQlt3npJm6NfwkaILVUygNOKheDIjxCBXNNzk5wFBl7yyFLcxdPNTnNipmoNbgDXEiJWQ9
3KxC0cEEskkRREKz/VtHLThoKuP4OK7EOavt4tdRQzByKi4DzfaDpcgR1q1hIfjv/ZM8uCzpwMaE
bhMllvK92D/1Jh0yM8CIYQfCpN03y7gO4GJ1Pp4PeVzxmFVojOjGBLkpM9U3dr97kvyQHcZbS/2R
o/ihFZzc2TaoSl44K90ucuP0u8Q2Mrt7z0kjgKY78HpGhaySCX7xodHkwfpsV5aYbmDIJ42moylV
Vvf/6beSWJs7QLSjCzMOitEgtlsqd8nrOfspdJNvY+MQvFsR32DR2k0rKJezUM4iUWuivKNXjk0O
DnMyvMDbPJR8+WFTYY1BTBNrzjFEdCMLrt+6sfWJ+UnJb8I6gz3CWxTBTnRfLQOnL0dcI21DlIxQ
cky1eDUzFtgWQHefwjwa5Vew5ZzpFFG/Cy9WdL3eoPYDdStUJUDOaJ9agohR+fvu39mkac7kjC8E
1818oTXUh10QZytimqshflZml/9IWxW5BXz6ZgxCadk9tf+cIbbFlUoDTUd5nSQlHmSZ4G/yhAVe
yd5jgz9dWnsIhioiWqk1Qze/nLr3sHUOsubS34O+ONC5YIUEeTUdX2rhXuNBS6EK8GFLdhnwVZPY
vuBlomxI22fs7yAeH9Dyra8xOC4NaJykF7QvPPaW8ohITYdx7YY6qgJfqyyAuKdDyYqkqc75EW1U
USzTyqXwReyfGzmYKFkc4eQm8Il1Dr+3JexjGvMTDhOtMJr078vqhv47/VchyqzbCWP8lyHRhpLH
ZXrY7JXiR+4/pFV6YhpMYF1F6XOw54z0wlS6rHJyX49iPYKR66tBMtoTruITn19z2TL4W9/HPGTT
imec5WzdvjSYTqfozVp2qcnXhot2j63EkD3X3TY/sl3WaX84Yt6jSzfs9A2rDSBgx1Jea08v8ZUf
ZUFfFJm5R9FATW3FqjzGu85dHWN3CNCwMJy62ryzw9zhxNaS+tz53lAplnRa2coBsSrljqEF+uO7
xJvv7qIZhNpXDGBfYzh+y9ACOGZy9psyeL4nrYpqozhi86d2HxplgO+a6A91tDVhXGSng4llI+CL
NqO5lCoIdS5A6IhSX6eh7MNzM6udO4pnCWk9MXbkG9NXNsvlzF4gdKy1n9YVMt3oFaNOYbq1y8Aj
1wcTvo5AjBdoejFMuXD+nupzKB2e+yyiXxybqVD7J/dphk8EWaQfdbt3XJ9/QPnPYZcRwj+ymezW
zzcyVuNYRiI+IG+nYzMELi6nJqDNUB5/rnK2dz1/XTGvz/G2RnjrplnF6EGt5/XiyhH0vTx9Bdum
3YUtQiLWD1sZwYW2eaDlA66qSdLgIsc/19L+OtZxsj+WeZylTJxNzjRt7XRjcC/UAMxvwWMUHBjd
zQFG8NWmNVkopQmmbZ7PQIWK33WJ7/Mgx+XwZftEsT/56iP0cfey3KRvfPZ7fdz5n35AgDWjO9yC
vZURNsGYg7ZJ40HZW7osCxaLo8/XYLMMjEAf1QsX6IRbZ1l3XLus5sfxnPp1S7SfiwRAPYyqRiVh
lL+bMI3Fu0fXzRcE3YTpVKOoJHoNQJ9p9P1Q1KfxwPF1JxJPw8hSODw5thrJqbpgWVSWM16BQ6LO
2Hbcbwdhg0P+frIAXPLthvv0YJ8D5lnQIXS3As878HmJ6+aQk6tSUNAie+D5+uaXjFIDO558qsJO
u5mqH/rnB/YuHxGvlLqFzTo/Hm7GLX5CQDVC+OUn1eoYbaAW7yOyh1nFumNZqSuSkcS7NYrexcCk
euHVY25Hz3ffWlUrM2Id/fNvbp8xEtuPZI4cD6ZZTAZk3w/IVZ4cF6IiDa2AX2eVADBIn01do7G7
Y4FK3zytX51b6PtxONGIss7bS0/jjZ6cWHMxWkBnIJjrOSItiqVyeVWm4KolgwRw2QGNFqmAHxhn
wV+Gxn3ZfNaILd8qPJIpIdKQ5hJVq+EsPLFW9/QAqEMlWFXbC4O6qA08OPO5iG2bal2FP5jlcTnD
3+10Q+zC8igCggI2KxbLWCYKtTzFg9KdDwGusoZvrOJxHVtTfRqc8opPshsf7SWKkKKdUl2LfWdD
cQb6yevfVRAZYdAersFzXsXXqtibBZkt6f747lOwVJO4s697gB6uKb6fGJbxV9uxlR+TohBXOGO9
JzD4xIc3pqWfogDaQbl4OTJyFM8a9AhvtQBPDD7741XUr7DtLDFunuvTr12x3tpFx/fio5OFR2EI
m/i6gWFXfU9uz+aiTikNFH213YKrNpPa1yYWq8jydrDJ/n8MHDr719m/MPHXnrqmACAqqGwJdUct
WvVlgZXiUBWRqoHvFRZsfrq7505rEsNoNbn8w97jK83bRZkfB2rUyQs2U6bQ4TUy18AnY0FWPwER
31xbuMHJ15tf7jkvK5RawlVlIRmhW2JaVVrgn9W55rgpxfYwt0Orq3XGW20RN1+1IEoFzWeaSRX5
ak1YW1rZTZ6CRRW8xEkWWknPaTdFs6BC48X+gRVoV85yMII6OFBrSGqY7CMLCWpMZs9A+cGoGDj9
ifOriwbiWgO1IR2536XYkA6B2fy3x7VvkS+/QppjBNQKdIRkWxgN9XiTJtr6BK2e2GpbhqiOzCgp
k4PXcCxIOMv5YBqXCfGObg3agVIcXu/TZXpTeb2cpsMddo+TOBrD02J8pBrKxcpFNNtcIrSRg9od
tGLZRxbuTWXJYpeT2qqT+6zFe44eByx1a/vquIAlxjBNAY1zZe4gAgOZRg7UpdtoZ7F82KAUu26D
wCYz2GXsgMmu/ez40y0SAkavYvbegv1VHpLvd59UAjW38BYBmLGKWHVzVuUUqYDUvLfE8/xnoAiS
RnOFqRXtlzEO3Y6GyCwOgDhwzPHpesMLQsAIz4DVR6I/DYq40pbz8ZfbFupiqwPOGD9yEQmcN8+F
ONPENfwdrz4LbpVWe9CqVElob+Gm+mnmhiCr8f7G6UYhH+AwwZBtym7KXVJ7Y/7h/oN9X4B1WMj5
cGUFhvsrYlSA/O/392KDEIF3FD1tQIALjePyl/REox49Kaesz9YrrpcpCXr/D5E5hUsR8U6fTkAE
JeBaTdr3VeuKylSkPpjyZsztpbHi5Gqxf9fYjIETSMt83ul6eCkZKvTbYN4DvbmIeJ8YSkSv+AcW
Lt+Oe1vajHdMp+uZ5W6r0zZVDao/6a8eNnl21D2S0AGzm9GxsnYMxuzVg4q2HEWpVZABd5E88PpX
jaFcnes0NMyjnEwIi+q1nQgKGa3yp3Wg7tvTAADbLsr3T22DQBVdckpv1UrF0iEEUwdF/Fe1kjKF
xUIN41dQ1pkytzHHEEZ2QwFA6u7bQI+LyWueAoGO0y8tUOfyNVy43Ux2QF3EgP6vXYUYIFqA8Z/7
FmDHDxYBykaPkh4KpH7pht+XJ9ZAoQz6HkQ0F5dEsuuhsdJbfzNbgnn0BJr+1wA7zwzILWCuEFaX
87nqmaNeegI2T+Ktx3YBXxlILvdJDYd3vNhJc7KguXdQXNmnftStx/h6WsjB9L03PpB93Rcv1ICi
PvdGeT/41RqcQrL+NypHKbk59Ny4NUSlKlfhZkDP1yOxFb6km7pkwYtBx71T+/yBRFbvr4y1WlPh
4JOn+1lr/7v+bA1VHKwuATvT8XXX1TDLjFdvp/2udZgjh9C2r3/478IePVyKcJ6GN0uLHWhdhbQ1
ItHA/EUsrETujlJ4/Q1nIxZ5zSaHdxV65t2mPFFWhtC7bQX2ogDRk+QmEr8W4m7rRYO3htSf68Dw
EMgpigcC/Cn6eqIaGYetpn9oMr8S3SYsw5k2+HsWD0WGWC3itYP3sfi2kQkVgiZDXWcYolc5KB7r
Oge+QpFkv2Lm/QRbOsp31UQpRS60Zoxt7iAn8gI17MYacqIBxxjJa4J8MzaxTMiPFGR1qv6rSlJq
NDtEVKcPdw5UR87xKGGMK4ZWzpT1z8vO+fZHQLOWoJZJHrCaOmDnQP6whlPZLnl181FkF81p2LMj
9A463tVcGwELApu4F8y2Crklyvi0cnmdLiRrtNjgTBo9HumenCJsvJ3CTXMcLec0/9MgPcG3X0T1
cjO4EcbrnjGmBQQccNOAp0R6fpedSYT4lJ5nC10INcTYx20wmLSxjGvhaGn/FTX7C4HOO5Q3FVHc
k72Rpj4DeCxQJC+44xTlT+IFqFotQCOagrhivu/UHO8cm6X4r9mE2tzoWRmvJlgGkANiD8Lq20jU
gDF6IYeg5+YZJIzMUKvFbqhJSz0ZegioEFZnHegy0uG/kt9YQzeVZuXEWn1YsBOr9WSsuHuaelyf
quwlXlyP0AJhrY/zztrLMuwoLwyD/taco7TVe/r89gGRSE6P0iNr9KYA4Wc4IrH5e6uln0pwgffG
BdmPbqutBQ2tJDvKNygJ+GLNciw+MCgYCOChYv1hOkNuTNzM7oyfYnhebTWjpCbpG+bpNlPVw/aw
yUyBN/mNgh9N0RLJztXstZ8eXSotWiPdn686vuHJK2reftV328CUotZaPBxFjA7m5Un+l+TQovus
YnxDqR+jSjDuSDrmyQMEQVK6Ttn+5/2Eqq6r7W8yyGyNkkXzUcnZMU+gdcJES+u5r5zmkw8SrJrX
ueLrtjbp7d1BGoCbi8Bvxzaee50yHc4g20Hx08BefyqIModGmaUHzPMw6k1+F5clbhrbREoPHCOp
zklGNTF8p7LMnp/RLDVC3r5cbS4NYrYLHEWh1R46rOd+MTLmq6rZ2bwlDGFO5W9Hy4LUOUMfRZk3
2FTWYB6JHh6QNGVGzyg4IPXdq/oHmYD8YnJ1YSy7CII59OeaPUbvkLZaxpsOSBFQrjhQiHxfHOK0
c7IZ0PkTLY2KtBphTtbE5GHkb3Su87W4g0y1oLnzIfNX3JVOCfqmAB64tKxI/iFSpfQuNwej2Qh7
FnCelcShpurUnuhzJHCsOKpe8OdSZkzFx64yJYEZN53KRdM+otMd0ThzBm3tC2B7eMbpL5E1ukKY
QjKfLGOaAb7xbI+MJhkynKvKqBBBJGK5xG5VD+Qlj2YRwU5qwbwnbhAXKEnP+brU3B5Lo3WwyWx0
MBmF0DG4NoN1RjGhE7+w839evYRPPRUK0ZpOJXsi8gqxDjTaO+eWpKzHfLWkocOMF38+/TRl/2Zo
p3vik7NXDHkiTkne1b7VbZ3M3Y0ifysrvSVV8/zs46y9PMtU68R0Goio/xbu5d9rQNYlc72IzkhG
tpjZ2MTZEMIhP5VavNgkkMssYgq3ngtDuBUx/IY9uHYKv/Lkqt/iRuYSE+6zPZMhdVyaCNtpGHlu
7ZmorXyeQQHBhzhfYjRC7uwtHJzz1Z3rKLmcAa1TPKrRSxGS3obhEr09TDM+jeB0NHkVdYMlygJU
Ip6uUhI6YL2gOpP71E4Alkr1mg3SQM3FcmVC2NxAuo2xujDzMde26CV2PPODQkYgMCTO7xxDbgHj
Ul2tPJNAHf8G6OQiKzj3rJxYLutamcxVDmKvA9tzz/FIDEWivuN8ZAaiUJC+7ffKCiV2v5wZXI2T
JZK6FEjdYoR/VkX1sSe71z7bMGpHdhfi1IKJUJ08+Q81BOqdLOH/QGvgDupR0V6qwvgMr5h/aZeW
XOk8AtxmUtrGjPBIT3GO/wjyhjWRYF6acxjL4EoC5yKzJua3rikbhXTykiNOGPQVOswBO+SvBcl3
sGAVRxJohrcwwTp5wVi4N3T6jrT8QJVHAde7xV66hAmWQvh0nfgCCDTJ22sunRpKojyWCLH8IT/D
yJ/Ie5vEcYgUciMVS2ewelRUtPLuVhk8nE52xwwxN1Mhsc1f55kkzvrvJn906Tot8FHFlNBtqPNg
eSTOAdgyd0sdRKYZh2cH+nfysIR/iI3HO58C70uJDpMKJeR7PnWMnIB+QBhP2gcOf8M2KQQ9CXmg
CPNmuVAXNV9WHChukaeAkm+wly4jJ/WVfub84gviRpTlhJ37AZv2MZRERTCVjWQuJJMk7UOr0OmG
s187OvKPHi6gwVRa68nGXLqgOjnTKyvEzCmQugt2vtbqhN/ddwRoMtrZF2v3yxbZmBlOF1u43dd4
iVOm4hfhI6rZrxMp0/PYr5x1ApJOqOVjITBE2NQLbBe+ULp0rSU5V5GTtgJJl84pVCRf36GUVo8C
Cf9O3LWeqNZNe1ICAVINKJF0s8H15gZLn16u1bS1reRsu9hb0EKYXpP0PSRWWMPSk4kN5V8Y739L
G6/ozAeVsHQEE/fcEyHWwFhSNGMY5/7jYX5DweZTUBicOCb0ni6zBPUnnSFfyydNpN/t17WK0Laz
YPBBxAmpGX61bnvA5A+KARjhozHTqd42IBQC1uOooiqhYTocHJ5KG3I/Pve2bn7ir88bjV2B/lSy
2a5ZMfYPocRWflrTthCnfk9btMk0auE/IwJ9Jt1CDdJ3g+DU9I9k8h9zR79+l+o3ER3vyQhZ8v/Y
6rwh40tmR9Ro9Vpa4CLt51Zw7fkVr/OZBs0bRUaNT9CZXsei397B1JGVimTQ57DtKQ0z9cPRJoPl
RmP/5GAvNuJMRAMfy8iBw7rDZa6JyjrEZcB6vupU29VorG19uqTJ+JA28zLoPIaDlHZ+RFTKfV1f
17L2gIifr8Ps3yEJu2yzZBQQdNVotbRYcHaBoui+np3RQ38A/4WqihFMmtxwWnjeFRTy/Felp7iS
4C88yJJXuSEL43qKtpD1eD5wb/4p+NVTMnmdYnV2VnFqdjYWkkYEGM8kcSiO8vjdAW41X+CaQNLF
i1OvHZ/OKAKuKZJaD9zg94E7sS38E3WnBeyLPoi77nzxTS963KEiKVJ32lXCKInwarCUyu1gQTdv
v/PFAZb/tSBtpSKsz7XfFVJD6RKhNtte9KEZxEZrfjoeusP/q+uwvHQ9G7QjWf/yG/cUfoMBMsG+
J8STtZA9YYtZOm0HexT8QvA0LizLYygcLeX6/na8A+B8D4I5KMYgIH5GWl53ALL+LSLKk9PAoldz
KSrHEnOs/+7LS/ef1NOYKDiZawCPp9fxk8nBrklvtFbKL/nwc4kVkQAbf2V+iNycx1fhMMqg7yzx
RlPuqUUXcxNQm6KJzMiz87/aVnDp6YW2rZnFNS5ORrG7mTDoZfRenmD6hjKd4h0hTBbRDqEm6jmW
BKsj4tU26RKdiRQP7bdDuTD/xwaa1CJdLOgTZ5/vZ9PqhMEIiRkiMdGdk5JPxrwy6M0hpP459ahn
G6V+lTitYBK2ulkDpsBMDq7/gIN1qamyGAIfKuQwsXQ2owvyXaLqBRBF+2y5m5DKRlzztohoH9kq
QREyFjOeS57Yk9GAVz91znyx4ho7YG6oTKhOxGAMH4F3IlPsLWCKt47GcrGw2Ygm2Kt62XPfrYtI
kFBc8SS4k8vm9TDo5gqdL1wMoFjNFd6sOi2CEAV7V6SfKlSAvuXw2jrKam+m4e1nRMXE6lRfrK33
u39khSmLvCDShNPuerAMlPYP+0ZDMB4vztvwMeoOv49rDXRLjEJZPyorav6335uZPJg0PAofPLCN
DNYCf4zwR6pugKPFoDKzNScp7sSD24gO/Il/bKVUWdKDtj+BRjB+NIxd534GwSVnfydNd5XnBlSu
/rZ0oM41r2WY1YaqvNI8L0mkGDTc2C5XvaMx+E1eeTwfsFtSwkPgy9fOASAoKZkYvMD8xISSOf9D
8N50y5rMY9V8Sm7A31eAmx4rfcJFVGdsFjqmvuWRgPVVGZuIMc1LVyFSFPKjNAO3j9KsmzJghgln
anX44x9B07Nf7Dpt+gkbIOVheNapw0tGXCXm9NHxh8IDG47fxFmccxnAd3lzLxPcSVIDU1mOz/MJ
JLPnDg5g+HNoBAeWJ+ykfnLpw1MlVqf2wEWojf/NRcOIOd+zF/1ub/AwaqPCRyZiahnTHus5T+HS
tQ38UbktPjcitbmfM25wlPg2R1lU/3QwHZ10d4oAltrb8miBE+LJfkgkOsUEeoVhljhYW87tUF/K
i8x/27mIXlUZQ14VGZHFK/8X+Nz80TPygJkQXy5CtFJvkma7OqVxGgWTQLLHi7OtXrCuCEQdmGQQ
ElnGOvWY99yGaIAGebmsvIpzc4auA0eqI3Llb8i+zNAQSQSnEqYq1O4N//i1YDP2HjWkPwaTmd/T
/vVxVMs7w4WQdHCp+v5XQRFn4vYPgwnxP3lD+b78Is5Gai/tN59QVZCIGkd/2+sAlYoWYmeaAqmo
tn11WyVxYeoxEOLyuFolPBfzXi0GSNWjD5mCcNEGzx0pdkZ5h7GGOYH4/QXfda0ZK3FvBj6WAu2I
wT/32wlzOtWOanW/otdjjQ7xIO0giPIcA9uWdDZa9KPj6+Yu/DJfG7PMevsti5iLgqXwQvy6Fp1E
Boc6f2YxpQfNOIU31XrhQ1Pn/gbYwYXwkHj3UNQEoznxF2Ipkk6ZbY4LZEHu/78DeEjTqxJZrt+Y
71NtMnbL39z505N1XdXB/XJEC3hKbgC1rsmeHfQVihw6aPU+XVpFxqU8k2ODzX/o5GIT6AE7vY1x
Ftj1rWx6QQRT7O2V/L5AbG6bYlVzVDhiys5c7M/B68XmHp9/HrRLN8qEIcPGmbNeub0L9vsKk1eV
iaOf+vNV5js9sodCmE0um/0aeTDLmGFvL9G0b+jTIXO4ieM/0KdnYryuYeonzfTMOOm6YyGqihfB
8Vm03AY13PgKyRq99Qh0TBJxbKZrCFNRvu3e+eX2wteus4CYQ1ILRZ9eHiSKEelUanY5NrxddeK5
JTV1kavtyTqM9jF9heRzmi4jb4ZewtNateT7tsdfcwipJERIN48yjhN7bcpX3MiCO805KyZenDd5
AAXc+8z51R42ng7UEW/rKOc6ilQPKWp9reAq66iCsmUHapPRs2DKAb0ax5Ok1N5yK2WLsT7Mu+ki
4Vcb0xjCCFD0W96cV1fhvzfblIJi8nGm4/XtbMFv94UbVh0OS1eJPbvI+IrV2Qg1fOj4v2D1my+f
nvPmqJrYVegM0jkcBr7J69nAlFRlzXwi2vg+NFQFgwG8xyEE0CeLTenDyTlUpxchMroP9OwfAUMp
2TjQY0QeJoV4B2hYa88AFqiRoeUOzwzSkVWqoYBbJfoBISmrTOSteEd4rY0EC8cbJRErYTiozNeQ
Hdad0drzvgSdkEo3yk+KcFdIpgU/MBXeYyCRifc3mSQULH7/u5ud8U2xB1aQ6Aum+W5fw4XHqpY5
BJSiM939mo4UPLyrkcSCAMcPkymmotLhzQ9+JZJblzE+ZAMmj0WPHzRJT/PmXKkjIhd3pvH2jkwY
oVIa4pcwukZmWPb4S2/OFI+8RSMhpfjZqr3m3NOYRja/JuDFh857EFfEMQB/wXbG9paWsI4wfBwQ
XM7+TkxPX5LI/xz4GSPqH/3AwaBJBoxlKppxPawnk/4dYfKx/9x6/5CL3MUH+1NypktmcLZawyah
S2gsU42lfkMylQxzsjCzD4P0IhxGd7jFaH/7uNtmOIQm5ib0G9e6gbkQkW/HjclRC0JpjykShaqQ
izK4WXPc1WTW6HALVlIgSFPrkTukCCDP/9ywVNBLdAN5kX6fEamV02nJTeiGaHj4C0iFo3+Ivl2s
T4zbE2NYD8lzalGRR0Ude/pLbCiJ6QWvEVpWkgOp4iLF5/O2Foo1ZOWQAztP+oud7lTcMBWsxOI2
84eBOXbkf9XRPxgvGwQY8MSArMZmEhZ7qnJfDXS2d0IADm8gAX1e0TXa0NcKTefJ2Uoo5Kj4LeeF
Rem2+lU0r6gHO9bZjIE+aife5ME3appEONHlctRi/Q1faxWmqNWH1KW2nxUvikgcWpf3JssmQcNA
WMuKqyEkVR5Q1u0lFPNAseotrg/tP7SraCxtI/W1HS1ilp5wEW78xhCrEWctXYgCd+rpecqGfeoF
8RAv2Ju9MotSYpBlhGaMs2W5AiuknzAi/v8ZyuPSr74LuUootyB6Vzz+FUiJffOXz0C3PoZ28o9S
M6Aormc8jvdRp07ZDMhmqa3A4plRITB492BfXAGC67MPyK8funv45jj9jSphlCNcgqFyhFjL+1De
eSgvbCDVhNQhxD2573pu0NsbCJSUd7iz1K9uwOKOQZFJ8gbC6QqoAy3YTxZarw+fPyeG+gp1O99M
LddfRovd8HNNPoVbFXONSxTev3XMWo02sYneXu6rU6xKHtyNHXttB/UjfYNSQ0RXKbTjIYrc05VF
FlN2htjKNlJNMb7Q1lRP4QUFbdJ1y5KCgcQB+bLNefAydO+bJJaB91PSLgca1pi2peaiyZFYdtv9
bPLNKxQZJpWaovPKuylQL44uXd7bet3OxyGnN/s3ydG6q+qDx7VWy2frDWfUID7NJOl+JFaVKWGy
voFY+lkNKLc768RZXWo8pDvK+q77cYNaF0CMT70WtstnK8KB04BWuQeSx29Yfx79wByuKUJkLppC
g+iMsksCA33ISbzJRBEaaWH0ZXNdi4c6NDAox2r0gwFjoJU7GYMXr8b8bcUYbeJqUKImwB27hmnV
FuIQunzsRXS2wjzuFKfAXyENUgXHl5rvaSsJSePrN5c0OSa24buuoAGvlXFjopu1cHntf81eYecT
cY+Nvx7oiE1tVA+T/scVGDwdVmHLW+TnJo4TfqK9AdV7j76tKujxSy2aicY7k/zHfeJlXigvRtaV
pLdOiEhD+aaFAvwzKrpvvVnWsvWP6/UYM62A8PfqQ9qeeLwUUucBsWBCAhmNjto+g/tn1R4ceyiL
Q5sEenHkufgwsaFFTJ6ZqGhF3YbvEAZqDGUIzXKJI1yZeuxNRy5AwgFIC6AlNVsZAdxhEWE3MSOR
rcW3LNOEoTrAttfuovO3OiBOdQpfXO+MfDmJuBf1yQEzLJOA+f38OPWlbammL/U241MOo0tBUaSZ
GzeOS5E8QMcL6OFDXtBaxsIO2xjjR3zrBaAWcLVVv/ihb0mkmm66bZfrXjWG6As0BJsZhTxKrkao
9THbAaK0s5XMJUqHjrqG/EJkZDuI5atg0GEIuUDIKobvd8G4cKqrA6IwakXo3o5laVrPOCIzzBAZ
vIQdJ00qKsx8jon3NuPd4onpCB7MN2taNq9p1wUseKmK9KSq081bEfSemeHnE4bvyeB54pp7F8Mn
PbBCFtJnIpAT1TPpxU1zUH4J2MQ4JJZlMmkvVZpvo2jok0ZEHVduNYo8sKfF9ta4F6KoHzW4OHv6
B5WOCz5P6PfwM9N9sjXRSabvLChzPy3z0BEdbVyC1/k+HQgVBJ0yVoE6VdPbOUU+SCp9OJlQZuam
jPxgp9Sup5/YLRHhGwuvYyEfkFZDcYUbKqd590Nh310nYQSx8qtg93xpPkT4HgijPjrd7s5RT868
YTYclg6l2EdPs4GD1zPeveriYB9SDvU6wVpwyue1irZ0Ez5heIM8TxURi9YMvFsO3tsm6jKdD+0t
KRo4adkixhCpB62bykUjVaf37gChj6NV+kgIOnIk1LDJ5b7p16luM7aADYLu/wuCwrdcZw7o+Z6u
Rz4CmdmQy7F2VRHsxBd/bQZw8JZ6hcx8Tqdk39t4fEZ62iufsEe7xIOfxso4+HjDs7nd649NlJrO
ZEwB0hmluMGSN22ejkY1SnUZqqhKBDVPTHxR+TqtDltGPBHzrMQ80JaP47d88B6j1WJsAtaC5Jxm
Z8qDMW5OJ47K+64aFGUmERA8TGrMY15W5MG/EWX4anaYEedX7Hr4oLGZ7N2VNwby6ZZBpVt2Q7Fp
v8uXk4I3S2P/2SATAx8n3lgsFBPLfAuFSRNCkaIGpIqJrC+soHLldm4+toj2yURRxhAbnBsLWzvW
eNj76FDCd4YE6TBPYKu/j0aQY/NwT9BVoqf/y/Y1ToUfDG3BvRyWyU2kEtO4kQe4fINUrAByhmC4
9yrjjX9NhQf4oN0F6MCXQ5Fjn8CzEYnTLqP4w1AS5B3RoPMUZq8oCftrtYZ9EdXqSJ1gx2IQjFQi
LgdpskV10gWgjJ0GW2ITV+Y2ArlF44t3xoKp80khjeT+Vxs6uLr2iypP1WGffe+PD1r8CyE6/Bdy
KGxZfb7dK7b9Fy5APowS2cV47azrRVAyUOUAuqGi2a0znZGH/5WwKtcOg4WXukjfajEh0LXWXvpq
4+u3E08fTs4nvpdkeOCdsd7/UWl3WFR5+tFa7S4oKIR/dXDqEMRGafXbBc+0HeRS+5LpN1KmkX5j
7Pk+ggRY3uca+lTLUZj6O96RljACvBiUhJrTv2qSEIk3ysrJ1o3MzgyIAUlgB2VxYPeBo6t248HG
TxGmhCf/XmGzOppRSX2sF81Ljdy5zrs4sWSILZ0dgWRL9ygXl4Pqn+D4D7A3pZvXTTvq3wxju2S4
uEsRIoLUCI+xjpe6jEb6x+LPYqW6a8H92Ga5+FDP0uc5ILpeFQNuXob7XU9jXCK9le9F3AVl+ubB
FUoK5T6ajaFmzft+l+JFJBKQKLotvurKPVf9LpqzM+ILXtZvGSs/6LntOWgWkX3WqKR5lwalskcO
Zgvy6BrX8SrE/VdygsxB7sB59AMsRthzItzs5R7bTM+0A8fcljA0HHr0J1XfK/e1Cb/A+KN6xKPl
/E+tacDox+lxknxBYptJQ9G6zm6YhccqlqyC/B1/WRZuXqokFxguF0EvyLwlaNweJC9n946Ma+nY
ljDNoiLBC84dS3cFtXRJeBPEJqu9IHaRruzCfzKTLaSzHsEaGSU+ixuc6XA707CFMs034zPvi8xL
9WjlNvfgUqEs5j+oVTxR8GQDNrq+odfHXxOI+hlo3O53rN5CddISVH/D/LB0Vc72uoBbFoZHk30V
u1EZRaiU/3g7nuC0HGC6VxfrLXCQuDa4UKQkVIGkdKxeWYj/KXV6A7FIM3i9ETpluFVBZLZCQWhs
yWv3dvZ0eNyRRyfJ056yOYrn+JUp3ZwDiWELtYMDupZHHFswJRgMTA6skH/XXNuaBgZWrwLYnDfW
ef56w8IWj5y+bu2IAICW8k0TrMWz7/z1Oa/3U+GONZk0cIjoTOx2l083mOVVF0h94f3F0E1mY7/J
SnwAeNt/i37wzlvQZB5aimEPXgRB10yLAqakZCLNCflDC14H7RBzVpyEegrxtO1f55n5B9TWnvCM
KnE/z9AISdoXJ+8N5llI3BOOWtSA9r9cN4W1JbeoEH2ebrgUE8Ra5akkOIbqW7M2B485WUJ1Ltau
eopqXod+vXbIW2getu9lyowe6m+w8ocx8A7aS5wD7v16d9rFZCfis43EsFmsbsclpcjceUuGKvoa
U/ZeSj6qmlnrNPsA2mb3iQq4kS+16RqH7ZyteeZfc6w1lN5Zsyovf4hHQNM3bq4TLS22CtFle0RM
F2XDZmD/Kh6hC9nA6kAPxP54dYwAWbJDKPjro52dPUMcq+8en/oIRFzVocWwKQcuyRaR54uQoGu8
AiKIv3rBt84Hht6809EMW1WW8mNaExA2OC1n7RG3suLlCllNR6jD50Q+JPsHT4VGyvRNTwZFOjVo
Hphn+1HlhDQbPOyJdsZ3Gx/N97aON4xfsKvaZHxImzyW0RGL0y3hnxmdfovNPvFxDK6T6WER0IgU
yh9mlla/IyZDc0pY2PfR0f9jlWaChddvcynf4moHaxkxXIc1i9WFyrQ0AkJR8wfAetvDuQQryk7i
B5f1aeuz
`pragma protect end_protected

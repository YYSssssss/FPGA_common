//Personality Parameters
localparam  MAJOR_VERSION ='h0;
localparam  MINOR_VERSION ='h0;
localparam  REVISION_NUM  ='h1;
localparam  DEBUG_REVISION='h0;
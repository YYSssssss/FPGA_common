

module  lut_sensor_36fps_ir(
    input       [10:0]  lut_index,
    output reg  [39:0]  lut_data
);


//=====================================================
//              signals declare
//=====================================================


//=====================================================
//              rtl body
//=====================================================

//always @*
//begin
//    case(lut_index)


///* 11'd1          :lut_data = {8'h90,16'h0010,16'hf100};
//11'd2          :lut_data = {8'h90,16'h0322,16'h3000};
//11'd3          :lut_data = {8'h90,16'h0332,16'hf000};
//11'd4          :lut_data = {8'h90,16'h0313,16'h4000};   //16'h8200
//11'd5          :lut_data = {8'h90,16'h0316,16'h1e00};
//11'd6          :lut_data = {8'h90,16'h0314,16'h0000};
//11'd7          :lut_data = {8'h90,16'h031d,16'h6400};
//11'd8          :lut_data = {8'h90,16'h044a,16'h4000};
//11'd9          :lut_data = {8'h90,16'h040b,16'h0700};
//11'd10         :lut_data = {8'h90,16'h042d,16'h1500};
//11'd11         :lut_data = {8'h90,16'h040d,16'h1e00};
//11'd12         :lut_data = {8'h90,16'h040e,16'h1e00};
//11'd13         :lut_data = {8'h90,16'h040f,16'h0000};
//11'd14         :lut_data = {8'h90,16'h0410,16'h0000};
//11'd15         :lut_data = {8'h90,16'h0411,16'h0100};
//11'd16         :lut_data = {8'h90,16'h0412,16'h0100};
//11'd17         :lut_data = {8'h90,16'h0333,16'h1b00};
//11'd18         :lut_data = {8'h90,16'h0413,16'h0200};
//11'd19         :lut_data = {8'h90,16'h0414,16'h0200};
//11'd20         :lut_data = {8'h90,16'h0415,16'h0300};
//11'd21         :lut_data = {8'h90,16'h0416,16'h0300};
//11'd22         :lut_data = {8'h90,16'h042d,16'h5500};
//11'd23         :lut_data = {8'h90,16'h042e,16'h0100};
//11'd24         :lut_data = {8'h90,16'h0320,16'h2400};
//11'd25         :lut_data = {8'h90,16'h0100,16'h2200};
//11'd26         :lut_data = {8'h90,16'h0100,16'h2300};
//11'd27         :lut_data = {8'h90,16'h0325,16'ha500};
//11'd28         :lut_data = {8'h90,16'h0313,16'h4200};
//11'd29         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd30         :lut_data = {8'h80,16'h0001,16'h0800};
//11'd31         :lut_data = {8'h80,16'h0002,16'h1300};
//11'd32         :lut_data = {8'h80,16'h0100,16'h6000};
//11'd33         :lut_data = {8'h80,16'h0101,16'h4a00};
//11'd34         :lut_data = {8'h80,16'h0007,16'h0700};
//11'd35         :lut_data = {8'h80,16'h02d4,16'ha700};
//11'd36         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd37         :lut_data = {8'h80,16'h02d3,16'h8400}; */


//11'd1          :lut_data = {8'h90,16'h0010,16'hf100};
//11'd2          :lut_data = {8'h90,16'h0322,16'h3000};
//11'd3          :lut_data = {8'h90,16'h0332,16'hf000};
//11'd4          :lut_data = {8'h90,16'h0313,16'h4000};   //16'h8200
//11'd5          :lut_data = {8'h90,16'h0316,16'h1e00};
//11'd6          :lut_data = {8'h90,16'h0314,16'h0000};
//11'd7          :lut_data = {8'h90,16'h031d,16'h6400};
//11'd8          :lut_data = {8'h90,16'h044a,16'h4000};
//11'd9          :lut_data = {8'h90,16'h040b,16'h0700};
//11'd10         :lut_data = {8'h90,16'h042d,16'h1500};
//11'd11         :lut_data = {8'h90,16'h040d,16'h1e00};
//11'd12         :lut_data = {8'h90,16'h040e,16'h1e00};
//11'd13         :lut_data = {8'h90,16'h040f,16'h0000};
//11'd14         :lut_data = {8'h90,16'h0410,16'h0000};
//11'd15         :lut_data = {8'h90,16'h0411,16'h0100};
//11'd16         :lut_data = {8'h90,16'h0412,16'h0100};
//11'd17         :lut_data = {8'h90,16'h0333,16'h1b00};
//11'd18         :lut_data = {8'h90,16'h0413,16'h0200};
//11'd19         :lut_data = {8'h90,16'h0414,16'h0200};
//11'd20         :lut_data = {8'h90,16'h0415,16'h0300};
//11'd21         :lut_data = {8'h90,16'h0416,16'h0300};
//11'd22         :lut_data = {8'h90,16'h042d,16'h5500};
//11'd23         :lut_data = {8'h90,16'h042e,16'h0100};
//11'd24         :lut_data = {8'h90,16'h0320,16'h2400};
//11'd25         :lut_data = {8'h90,16'h0100,16'h2200};
//11'd26         :lut_data = {8'h90,16'h0100,16'h2300};
//11'd27         :lut_data = {8'h90,16'h0325,16'ha500};
//11'd28         :lut_data = {8'h90,16'h0313,16'h4200};
//11'd29         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd30         :lut_data = {8'h80,16'h0001,16'h0800};
//11'd31         :lut_data = {8'h80,16'h0002,16'h1300};
//11'd32         :lut_data = {8'h80,16'h0100,16'h6000};
//11'd33         :lut_data = {8'h80,16'h0101,16'h4a00};
//11'd34         :lut_data = {8'h80,16'h0007,16'h0700};
//11'd35         :lut_data = {8'h80,16'h02d4,16'ha700};
//11'd36         :lut_data = {8'h80,16'h02d6,16'h9400};

////11'd37         :lut_data = {8'h90,16'h03e0,16'h0000};
////11'd38         :lut_data = {8'h90,16'h03e2,16'h0000};
////11'd39         :lut_data = {8'h90,16'h03e7,16'h0c00};
////11'd40         :lut_data = {8'h90,16'h03e6,16'hb700};
////11'd41         :lut_data = {8'h90,16'h03e5,16'h3600};
////11'd42         :lut_data = {8'h90,16'h03ef,16'hc000};
////11'd43         :lut_data = {8'h90,16'h03f1,16'h4000};
////11'd44         :lut_data = {8'h00,16'h0000,16'hff00};
////11'd45         :lut_data = {8'h80,16'h02d3,16'h8400};

//11'd37         :lut_data = {8'h00,16'h0000,16'hff00};

//11'd38         :lut_data = {8'h90,16'h02cb,16'h9300};
//11'd39         :lut_data = {8'h80,16'h02d8,16'h0900};
//11'd40         :lut_data = {8'h80,16'h02c3,16'h0800};


//11'd41         :lut_data = {8'h80,16'h02d3,16'h8400};

////debug
//11'd42         :lut_data = {8'h80,16'h0001,16'h0800};
//11'd43         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd44         :lut_data = {8'h80,16'h0002,16'h1300};
//11'd45         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd46         :lut_data = {8'h80,16'h0100,16'h6000};
//11'd47         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd48         :lut_data = {8'h80,16'h0101,16'h4a00};
//11'd49         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd50         :lut_data = {8'h80,16'h0007,16'h0700};
//11'd51         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd52         :lut_data = {8'h80,16'h02d4,16'ha700};
//11'd53         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd54         :lut_data = {8'h80,16'h02d6,16'h9400};
//11'd55         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd56         :lut_data = {8'h80,16'h02d8,16'h0900};
//11'd57         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd58         :lut_data = {8'h80,16'h02c3,16'h0800};
//11'd59         :lut_data = {8'h00,16'h0000,16'hff00};
//11'd60         :lut_data = {8'h80,16'h02d3,16'h8400};

//        default :lut_data = {16'hff,16'hffff,16'hffff00};								   
								   
								   
//    endcase 								   
//end         




always @*
begin
    case(lut_index)
    
11'd1          :lut_data = {8'h90,16'h0010,16'hf100};
11'd2          :lut_data = {8'h90,16'h0322,16'h3000};
11'd3          :lut_data = {8'h90,16'h0332,16'hf000};
11'd4          :lut_data = {8'h90,16'h0313,16'h4000};   //16'h8200
11'd5          :lut_data = {8'h90,16'h0316,16'h1e00};
11'd6          :lut_data = {8'h90,16'h0314,16'h0000};
11'd7          :lut_data = {8'h90,16'h031d,16'h6400};
11'd8          :lut_data = {8'h90,16'h044a,16'h4000};
11'd9          :lut_data = {8'h90,16'h040b,16'h0700};
11'd10         :lut_data = {8'h90,16'h042d,16'h1500};
11'd11         :lut_data = {8'h90,16'h040d,16'h1e00};
11'd12         :lut_data = {8'h90,16'h040e,16'h1e00};
11'd13         :lut_data = {8'h90,16'h040f,16'h0000};
11'd14         :lut_data = {8'h90,16'h0410,16'h0000};
11'd15         :lut_data = {8'h90,16'h0411,16'h0100};
11'd16         :lut_data = {8'h90,16'h0412,16'h0100};
11'd17         :lut_data = {8'h90,16'h0333,16'h1b00};
11'd18         :lut_data = {8'h90,16'h0413,16'h0200};
11'd19         :lut_data = {8'h90,16'h0414,16'h0200};
11'd20         :lut_data = {8'h90,16'h0415,16'h0300};
11'd21         :lut_data = {8'h90,16'h0416,16'h0300};
11'd22         :lut_data = {8'h90,16'h042d,16'h5500};
11'd23         :lut_data = {8'h90,16'h042e,16'h0100};
11'd24         :lut_data = {8'h90,16'h0320,16'h2400};
11'd25         :lut_data = {8'h90,16'h0100,16'h2200};
11'd26         :lut_data = {8'h90,16'h0100,16'h2300};
11'd27         :lut_data = {8'h90,16'h0325,16'ha500};
11'd28         :lut_data = {8'h90,16'h0313,16'h4200};
11'd29         :lut_data = {8'h00,16'h0000,16'hff00};
11'd30         :lut_data = {8'h80,16'h0001,16'h0800};
11'd31         :lut_data = {8'h80,16'h0002,16'h1300};
11'd32         :lut_data = {8'h80,16'h0100,16'h6000};
11'd33         :lut_data = {8'h80,16'h0101,16'h4a00};
11'd34         :lut_data = {8'h80,16'h0007,16'h0700};
11'd35         :lut_data = {8'h80,16'h02d4,16'ha700};
11'd36         :lut_data = {8'h80,16'h02d6,16'h9400};

11'd37         :lut_data = {8'h00,16'h0000,16'hff00};

11'd38         :lut_data = {8'h90,16'h02cb,16'h9300};
11'd39         :lut_data = {8'h80,16'h02d8,16'h0900};
11'd40         :lut_data = {8'h80,16'h02c3,16'h0800};

11'd41         :lut_data = {8'h80,16'h02d3,16'h8400};

//debug
11'd42         :lut_data = {8'h80,16'h0001,16'h0800};
11'd43         :lut_data = {8'h00,16'h0000,16'hff00};
11'd44         :lut_data = {8'h80,16'h0002,16'h1300};
11'd45         :lut_data = {8'h00,16'h0000,16'hff00};
11'd46         :lut_data = {8'h80,16'h0100,16'h6000};
11'd47         :lut_data = {8'h00,16'h0000,16'hff00};
11'd48         :lut_data = {8'h80,16'h0101,16'h4a00};
11'd49         :lut_data = {8'h00,16'h0000,16'hff00};
11'd50         :lut_data = {8'h80,16'h0007,16'h0700};
11'd51         :lut_data = {8'h00,16'h0000,16'hff00};
11'd52         :lut_data = {8'h80,16'h02d4,16'ha700};
11'd53         :lut_data = {8'h00,16'h0000,16'hff00};
11'd54         :lut_data = {8'h80,16'h02d6,16'h9400};
11'd55         :lut_data = {8'h00,16'h0000,16'hff00};
11'd56         :lut_data = {8'h80,16'h02d8,16'h0900};
11'd57         :lut_data = {8'h00,16'h0000,16'hff00};
11'd58         :lut_data = {8'h80,16'h02c3,16'h0800};
11'd59         :lut_data = {8'h00,16'h0000,16'hff00};
11'd60         :lut_data = {8'h80,16'h02d3,16'h8400};

    default :lut_data = {16'hff,16'hffff,16'hffff00};							   
    endcase 								   
end         

            
endmodule   
            
module jb_interface_map_top(
    input                               syn_data_dl_ul_5ms,
	input                               tuser_dl_frm_mrkr_10ms,
    jb_dl_dfe_ctrl_if.dl_dfe            IFP_dl_dfe_ctrl,
    jb_ul_dfe_ctrl_if.ul_dfe            IFP_ul_dfe_ctrl,		
	jb_cmn_ctrl_if.cmd_dfe              IFP_cmn_ctrl,
	jb_oran_lphy_ctrl_if.lphy           IFP_oran_lphy_ctrl,            
	
	jb_dl_dfe_ctrl_devided_if.ctrl      IFP_dl_dfe_ctrl_new[1:0],
	jb_ul_dfe_ctrl_devided_if.ctrl      IFP_ul_dfe_ctrl_new[1:0],  	
	jb_cmn_ctrl_devided_if.ctrl         IFP_cmn_ctrl_new[1:0],
	jb_oran_lphy_ctrl_devided_if.ctrl   IFP_oran_lphy_ctrl_new[1:0],
	
    jb_axi4_stream_if.slave             IFP_dpd_s_axis_din[1:0],    // 128,32
    jb_axi4_stream_if.master            IFP_dpd_m_axis_dout[1:0],   // 128,32
	
    jb_axi4_stream_if.master            IFP_dpd_s_axis_din_new,     // 256,64
    jb_axi4_stream_if.slave             IFP_dpd_m_axis_dout_new,    // 256,64
									    
    jb_axi4_stream_if.slave             IFP_cfr_s_axis_din[1:0],    // 128,1
    jb_axi4_stream_if.master            IFP_cfr_m_axis_dout[1:0],   // 128,1
									    
    jb_axi4_stream_if.master            IFP_cfr_s_axis_din_new,     // 256,1
    jb_axi4_stream_if.slave             IFP_cfr_m_axis_dout_new     // 256,1
	
	);
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[0][0]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[0][0];
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[1][0]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[1][0];
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[0][1]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[0][1];
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[1][1]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[1][1];
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[0][2]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[0][2];
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[1][2]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[1][2];
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[0][3]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[0][3];
    assign IFP_dl_dfe_ctrl_new[0].dl_dfe_mute_path[1][3]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path0to3[1][3];		
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_int_frac_delay_trig             = IFP_dl_dfe_ctrl.dl_ant_int_frac_delay_trig;
	assign IFP_dl_dfe_ctrl_new[0].dl_car_nco_lsb[0][31:0]                = IFP_dl_dfe_ctrl.dl_car_nco_lsb[0][31:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_car_nco_lsb[1][31:0]                = IFP_dl_dfe_ctrl.dl_car_nco_lsb[1][31:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_car_nco_msb[0][6:0]                 = IFP_dl_dfe_ctrl.dl_car_nco_msb[0][6:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_car_nco_msb[1][6:0]                 = IFP_dl_dfe_ctrl.dl_car_nco_msb[1][6:0];			
	assign IFP_dl_dfe_ctrl_new[0].dl_car_nco_msb[0][7]                   = IFP_dl_dfe_ctrl.dl_car_nco_sign[0];		
	assign IFP_dl_dfe_ctrl_new[0].dl_car_nco_msb[1][7]                   = IFP_dl_dfe_ctrl.dl_car_nco_sign[1];		
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler_sign[0][3:0]     = IFP_dl_dfe_ctrl.dl_stream_gain_scaler_sign[0][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler_sign[1][3:0]     = IFP_dl_dfe_ctrl.dl_stream_gain_scaler_sign[1][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[0][0][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][0][3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[0][1][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][1][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[0][2][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][2][3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[0][3][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][3][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[1][0][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][0][3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[1][1][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][1][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[1][2][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][2][3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_scaler[1][3][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][3][3:0];																	     
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[0][0][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][0][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[0][1][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][1][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[0][2][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][2][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[0][3][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][3][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[1][0][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][0][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[1][1][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][1][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[1][2][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][2][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_stream_gain_fraction[1][3][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][3][15:0];		
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_scaler_sign[3:0]    = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler_sign[3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_scaler[0][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[0][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_scaler[1][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[1][3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_scaler[2][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[2][3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_scaler[3][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[3][3:0];		
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_fraction[0][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[0][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_fraction[1][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[1][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_fraction[2][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[2][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_precfr_gain_fraction[3][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[3][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_scaler_sign[3:0]   = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler_sign[3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_scaler[0][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[0][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_scaler[1][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[1][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_scaler[2][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[2][3:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_scaler[3][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[3][3:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_fraction[0][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[0][15:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_fraction[1][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[1][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_fraction[2][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[2][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_postcfr_gain_fraction[3][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[3][15:0];		
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_delay[0][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[0][5:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_delay[1][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[1][5:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_delay[2][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[2][5:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_ant_delay[3][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[3][5:0];	
	assign IFP_dl_dfe_ctrl_new[0].bypass_dpd                             = IFP_dl_dfe_ctrl.bypass_dpd;	
	assign IFP_dl_dfe_ctrl_new[0].bypass_cfr                             = IFP_dl_dfe_ctrl.bypass_cfr;
	assign IFP_dl_dfe_ctrl_new[0].override_postcfr                       = IFP_dl_dfe_ctrl.override_postcfr;
	assign IFP_dl_dfe_ctrl_new[0].ps_filter_bypass                       = IFP_dl_dfe_ctrl.ps_filter_bypass;
	assign IFP_dl_dfe_ctrl_new[0].dl_dfe_path_dbg_sel[2:0]               = IFP_dl_dfe_ctrl.dl_dfe_path_dbg_sel[2:0];	
	assign IFP_dl_dfe_ctrl_new[0].clear_sat_flags                        = IFP_dl_dfe_ctrl.clear_sat_flags;	
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[0][0][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][0][6:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[0][1][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][1][6:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[0][2][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][2][6:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[0][3][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][3][6:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[1][0][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][0][6:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[1][1][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][1][6:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[1][2][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][2][6:0];
	assign IFP_dl_dfe_ctrl_new[0].dl_int_delay[1][3][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][3][6:0];																	     
	assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[0][0][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][0][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[0][1][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][1][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[0][2][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][2][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[0][3][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][3][15:0];	
    assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[1][0][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][0][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[1][1][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][1][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[1][2][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][2][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].dl_frac_delay[1][3][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][3][15:0];	
	assign IFP_dl_dfe_ctrl_new[0].pl_debug                               = IFP_dl_dfe_ctrl.pl_debug;

    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[0][0]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[0][0];
    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[1][0]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[1][0];
    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[0][1]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[0][1];
    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[1][1]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[1][1];
    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[0][2]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[0][2];
    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[1][2]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[1][2];
    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[0][3]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[0][3];
    assign IFP_dl_dfe_ctrl_new[1].dl_dfe_mute_path[1][3]                 = IFP_dl_dfe_ctrl.dl_dfe_mute_path4to7[1][3];		
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_int_frac_delay_trig             = IFP_dl_dfe_ctrl.dl_ant_int_frac_delay_trig;
	assign IFP_dl_dfe_ctrl_new[1].dl_car_nco_lsb[0][31:0]              	 = IFP_dl_dfe_ctrl.dl_car_nco_lsb[0][31:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_car_nco_lsb[1][31:0]                = IFP_dl_dfe_ctrl.dl_car_nco_lsb[1][31:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_car_nco_msb[0][6:0]                 = IFP_dl_dfe_ctrl.dl_car_nco_msb[0][6:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_car_nco_msb[1][6:0]                 = IFP_dl_dfe_ctrl.dl_car_nco_msb[1][6:0];		
	assign IFP_dl_dfe_ctrl_new[1].dl_car_nco_msb[0][7]                   = IFP_dl_dfe_ctrl.dl_car_nco_sign[0];		
	assign IFP_dl_dfe_ctrl_new[1].dl_car_nco_msb[1][7]                   = IFP_dl_dfe_ctrl.dl_car_nco_sign[1];		
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler_sign[0][3:0]     = IFP_dl_dfe_ctrl.dl_stream_gain_scaler_sign[0][7:4];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler_sign[1][3:0]     = IFP_dl_dfe_ctrl.dl_stream_gain_scaler_sign[1][7:4];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[0][0][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][4][3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[0][1][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][5][3:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[0][2][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][6][3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[0][3][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[0][7][3:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[1][0][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][4][3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[1][1][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][5][3:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[1][2][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][6][3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_scaler[1][3][3:0]       = IFP_dl_dfe_ctrl.dl_stream_gain_scaler[1][7][3:0];																	     
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[0][0][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][4][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[0][1][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][5][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[0][2][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][6][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[0][3][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[0][7][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[1][0][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][4][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[1][1][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][5][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[1][2][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][6][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_stream_gain_fraction[1][3][15:0]    = IFP_dl_dfe_ctrl.dl_stream_gain_fraction[1][7][15:0];		
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_scaler_sign[3:0]    = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler_sign[3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_scaler[0][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[4][3:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_scaler[1][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[5][3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_scaler[2][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[6][3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_scaler[3][3:0]      = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_scaler[7][3:0];		
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_fraction[0][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[4][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_fraction[1][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[5][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_fraction[2][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[6][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_precfr_gain_fraction[3][15:0]   = IFP_dl_dfe_ctrl.dl_ant_precfr_gain_fraction[7][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_scaler_sign[3:0]   = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler_sign[3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_scaler[0][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[4][3:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_scaler[1][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[5][3:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_scaler[2][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[6][3:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_scaler[3][3:0]     = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_scaler[7][3:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_fraction[0][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[4][15:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_fraction[1][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[5][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_fraction[2][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[6][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_postcfr_gain_fraction[3][15:0]  = IFP_dl_dfe_ctrl.dl_ant_postcfr_gain_fraction[7][15:0];		
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_delay[0][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[4][5:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_delay[1][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[5][5:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_delay[2][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[6][5:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_ant_delay[3][5:0]                   = IFP_dl_dfe_ctrl.dl_ant_delay[7][5:0];	
	assign IFP_dl_dfe_ctrl_new[1].bypass_dpd                             = IFP_dl_dfe_ctrl.bypass_dpd;	
	assign IFP_dl_dfe_ctrl_new[1].bypass_cfr                             = IFP_dl_dfe_ctrl.bypass_cfr;
	assign IFP_dl_dfe_ctrl_new[1].override_postcfr                       = IFP_dl_dfe_ctrl.override_postcfr;
	assign IFP_dl_dfe_ctrl_new[1].ps_filter_bypass                       = IFP_dl_dfe_ctrl.ps_filter_bypass;
	assign IFP_dl_dfe_ctrl_new[1].dl_dfe_path_dbg_sel[2:0]               = IFP_dl_dfe_ctrl.dl_dfe_path_dbg_sel[2:0];	
	assign IFP_dl_dfe_ctrl_new[1].clear_sat_flags                        = IFP_dl_dfe_ctrl.clear_sat_flags;	
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[0][0][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][4][6:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[0][1][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][5][6:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[0][2][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][6][6:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[0][3][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[0][7][6:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[1][0][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][4][6:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[1][1][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][5][6:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[1][2][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][6][6:0];
	assign IFP_dl_dfe_ctrl_new[1].dl_int_delay[1][3][6:0]                = IFP_dl_dfe_ctrl.dl_int_delay[1][7][6:0];																	     
	assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[0][0][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][4][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[0][1][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][5][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[0][2][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][6][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[0][3][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[0][7][15:0];	
    assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[1][0][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][4][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[1][1][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][5][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[1][2][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][6][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].dl_frac_delay[1][3][15:0]              = IFP_dl_dfe_ctrl.dl_frac_delay[1][7][15:0];	
	assign IFP_dl_dfe_ctrl_new[1].pl_debug                               = IFP_dl_dfe_ctrl.pl_debug;

	
	assign IFP_cmn_ctrl_new[0].hw_id                                     = IFP_cmn_ctrl.hw_id;
	assign IFP_cmn_ctrl_new[0].soft_reset                                = IFP_cmn_ctrl.soft_reset;
	assign IFP_cmn_ctrl_new[0].dl_stream_en[0][3:0]                      = IFP_cmn_ctrl.dl_stream_en[0][3:0];	
    assign IFP_cmn_ctrl_new[0].dl_stream_en[1][3:0]                      = IFP_cmn_ctrl.dl_stream_en[1][3:0];	
	assign IFP_cmn_ctrl_new[0].dl_car_bw                                 = IFP_cmn_ctrl.dl_car_bw;
	assign IFP_cmn_ctrl_new[0].ul_stream_en[0][3:0]                      = IFP_cmn_ctrl.ul_stream_en[0][3:0];	
	assign IFP_cmn_ctrl_new[0].ul_stream_en[1][3:0]                      = IFP_cmn_ctrl.ul_stream_en[1][3:0];	
	assign IFP_cmn_ctrl_new[0].ul_car_bw                                 = IFP_cmn_ctrl.ul_car_bw;
	assign IFP_cmn_ctrl_new[0].frm_mrkr_gen_enable[0]                    = IFP_cmn_ctrl.frm_mrkr_gen_enable[0];
	assign IFP_cmn_ctrl_new[0].frm_mrkr_gen_enable[1]                    = IFP_cmn_ctrl.frm_mrkr_gen_enable[1];
	assign IFP_cmn_ctrl_new[0].frm_mrkr_gen_trigger[0]                   = IFP_cmn_ctrl.frm_mrkr_gen_trigger[0];
	assign IFP_cmn_ctrl_new[0].frm_mrkr_gen_trigger[1]                   = IFP_cmn_ctrl.frm_mrkr_gen_trigger[1];
    assign IFP_cmn_ctrl_new[0].dl_frm_mrkr_cntr_ns[0][31:0]              = IFP_cmn_ctrl.dl_frm_mrkr_cntr_ns[0][31:0];
    assign IFP_cmn_ctrl_new[0].dl_frm_mrkr_cntr_ns[1][31:0]              = IFP_cmn_ctrl.dl_frm_mrkr_cntr_ns[1][31:0];
    assign IFP_cmn_ctrl_new[0].ul_frm_mrkr_cntr_ns[0][31:0]              = IFP_cmn_ctrl.ul_frm_mrkr_cntr_ns[0][31:0];
    assign IFP_cmn_ctrl_new[0].ul_frm_mrkr_cntr_ns[1][31:0]              = IFP_cmn_ctrl.ul_frm_mrkr_cntr_ns[1][31:0];
    assign IFP_cmn_ctrl_new[0].prach_frm_mrkr_cntr_ns[0][31:0]           = IFP_cmn_ctrl.prach_frm_mrkr_cntr_ns[0][31:0];
    assign IFP_cmn_ctrl_new[0].prach_frm_mrkr_cntr_ns[1][31:0]           = IFP_cmn_ctrl.prach_frm_mrkr_cntr_ns[1][31:0];
																	     
	assign IFP_cmn_ctrl_new[1].hw_id                                     = IFP_cmn_ctrl.hw_id;
	assign IFP_cmn_ctrl_new[1].soft_reset                                = IFP_cmn_ctrl.soft_reset;
	assign IFP_cmn_ctrl_new[1].dl_stream_en[0][3:0]                      = IFP_cmn_ctrl.dl_stream_en[0][7:4];
	assign IFP_cmn_ctrl_new[1].dl_stream_en[1][3:0]                      = IFP_cmn_ctrl.dl_stream_en[1][7:4];		
	assign IFP_cmn_ctrl_new[1].dl_car_bw                                 = IFP_cmn_ctrl.dl_car_bw;
	assign IFP_cmn_ctrl_new[1].ul_stream_en[0][3:0]                      = IFP_cmn_ctrl.ul_stream_en[0][7:4];
	assign IFP_cmn_ctrl_new[1].ul_stream_en[1][3:0]                      = IFP_cmn_ctrl.ul_stream_en[1][7:4];		
	assign IFP_cmn_ctrl_new[1].ul_car_bw                                 = IFP_cmn_ctrl.ul_car_bw;	
	assign IFP_cmn_ctrl_new[1].frm_mrkr_gen_enable[0]                    = IFP_cmn_ctrl.frm_mrkr_gen_enable[0];
	assign IFP_cmn_ctrl_new[1].frm_mrkr_gen_enable[1]                    = IFP_cmn_ctrl.frm_mrkr_gen_enable[1];
	assign IFP_cmn_ctrl_new[1].frm_mrkr_gen_trigger[0]                   = IFP_cmn_ctrl.frm_mrkr_gen_trigger[0];
	assign IFP_cmn_ctrl_new[1].frm_mrkr_gen_trigger[1]                   = IFP_cmn_ctrl.frm_mrkr_gen_trigger[1];	
    assign IFP_cmn_ctrl_new[1].dl_frm_mrkr_cntr_ns[0][31:0]              = IFP_cmn_ctrl.dl_frm_mrkr_cntr_ns[0][31:0];
    assign IFP_cmn_ctrl_new[1].dl_frm_mrkr_cntr_ns[1][31:0]              = IFP_cmn_ctrl.dl_frm_mrkr_cntr_ns[1][31:0];
    assign IFP_cmn_ctrl_new[1].ul_frm_mrkr_cntr_ns[0][31:0]              = IFP_cmn_ctrl.ul_frm_mrkr_cntr_ns[0][31:0];
    assign IFP_cmn_ctrl_new[1].ul_frm_mrkr_cntr_ns[1][31:0]              = IFP_cmn_ctrl.ul_frm_mrkr_cntr_ns[1][31:0];
    assign IFP_cmn_ctrl_new[1].prach_frm_mrkr_cntr_ns[0][31:0]           = IFP_cmn_ctrl.prach_frm_mrkr_cntr_ns[0][31:0];
    assign IFP_cmn_ctrl_new[1].prach_frm_mrkr_cntr_ns[1][31:0]           = IFP_cmn_ctrl.prach_frm_mrkr_cntr_ns[1][31:0];

	
    assign IFP_oran_lphy_ctrl_new[0].dl_swap_ifft                        = IFP_oran_lphy_ctrl.dl_swap_ifft;
    assign IFP_oran_lphy_ctrl_new[0].ul_swap_fft                         = IFP_oran_lphy_ctrl.ul_swap_fft;
    assign IFP_oran_lphy_ctrl_new[0].prach_swap_fft                      = IFP_oran_lphy_ctrl.prach_swap_fft;
    assign IFP_oran_lphy_ctrl_new[0].dl_iq_endianness                    = IFP_oran_lphy_ctrl.dl_iq_endianness;
    assign IFP_oran_lphy_ctrl_new[0].ul_iq_endianness                    = IFP_oran_lphy_ctrl.ul_iq_endianness;
    assign IFP_oran_lphy_ctrl_new[0].prach_iq_endianness                 = IFP_oran_lphy_ctrl.prach_iq_endianness;
    assign IFP_oran_lphy_ctrl_new[0].dl_ifft_gain_override[0]            = IFP_oran_lphy_ctrl.dl_ifft_gain_override[0];
    assign IFP_oran_lphy_ctrl_new[0].dl_ifft_gain_override[1]            = IFP_oran_lphy_ctrl.dl_ifft_gain_override[1];	
    assign IFP_oran_lphy_ctrl_new[0].ul_fft_gain_override[0]             = IFP_oran_lphy_ctrl.ul_fft_gain_override[0];
    assign IFP_oran_lphy_ctrl_new[0].ul_fft_gain_override[1]             = IFP_oran_lphy_ctrl.ul_fft_gain_override[1];
    assign IFP_oran_lphy_ctrl_new[0].dl_route_c0_to_c1                   = IFP_oran_lphy_ctrl.dl_route_c0_to_c1;
    assign IFP_oran_lphy_ctrl_new[0].dl_lte_5g[0]                        = IFP_oran_lphy_ctrl.dl_lte_5g[0];
	assign IFP_oran_lphy_ctrl_new[0].dl_lte_5g[1]                        = IFP_oran_lphy_ctrl.dl_lte_5g[1];
    assign IFP_oran_lphy_ctrl_new[0].dl_extended_cp[0]                   = IFP_oran_lphy_ctrl.dl_extended_cp[0];
	assign IFP_oran_lphy_ctrl_new[0].dl_extended_cp[1]                   = IFP_oran_lphy_ctrl.dl_extended_cp[1];
    assign IFP_oran_lphy_ctrl_new[0].dl_cc_numerology[0][3:0]            = IFP_oran_lphy_ctrl.dl_cc_numerology[0][3:0];
	assign IFP_oran_lphy_ctrl_new[0].dl_cc_numerology[1][3:0]            = IFP_oran_lphy_ctrl.dl_cc_numerology[1][3:0];	
    assign IFP_oran_lphy_ctrl_new[0].dl_ifft_scaler_sign[0]              = IFP_oran_lphy_ctrl.dl_ifft_scaler_sign[0];
	assign IFP_oran_lphy_ctrl_new[0].dl_ifft_scaler_sign[1]              = IFP_oran_lphy_ctrl.dl_ifft_scaler_sign[1];	
    assign IFP_oran_lphy_ctrl_new[0].dl_ifft_scaler[0][3:0]              = IFP_oran_lphy_ctrl.dl_ifft_scaler[0][3:0];
	assign IFP_oran_lphy_ctrl_new[0].dl_ifft_scaler[1][3:0]              = IFP_oran_lphy_ctrl.dl_ifft_scaler[1][3:0];		
    assign IFP_oran_lphy_ctrl_new[0].dl_ifft_fraction_gain[0][15:0]      = IFP_oran_lphy_ctrl.dl_ifft_fraction_gain[0][15:0];
	assign IFP_oran_lphy_ctrl_new[0].dl_ifft_fraction_gain[1][15:0]      = IFP_oran_lphy_ctrl.dl_ifft_fraction_gain[1][15:0];	
    assign IFP_oran_lphy_ctrl_new[0].ul_lte_5g[0]                        = IFP_oran_lphy_ctrl.ul_lte_5g[0];
	assign IFP_oran_lphy_ctrl_new[0].ul_lte_5g[1]                        = IFP_oran_lphy_ctrl.ul_lte_5g[1];
    assign IFP_oran_lphy_ctrl_new[0].ul_extended_cp[0]                   = IFP_oran_lphy_ctrl.ul_extended_cp[0];
	assign IFP_oran_lphy_ctrl_new[0].ul_extended_cp[1]                   = IFP_oran_lphy_ctrl.ul_extended_cp[1];
    assign IFP_oran_lphy_ctrl_new[0].ul_cc_numerology[0][3:0]            = IFP_oran_lphy_ctrl.ul_cc_numerology[0][3:0];
	assign IFP_oran_lphy_ctrl_new[0].ul_cc_numerology[1][3:0]            = IFP_oran_lphy_ctrl.ul_cc_numerology[1][3:0];
    assign IFP_oran_lphy_ctrl_new[0].ul_fft_scaler_sign[0]               = IFP_oran_lphy_ctrl.ul_fft_scaler_sign[0];
	assign IFP_oran_lphy_ctrl_new[0].ul_fft_scaler_sign[1]               = IFP_oran_lphy_ctrl.ul_fft_scaler_sign[1];
    assign IFP_oran_lphy_ctrl_new[0].ul_fft_scaler[0][3:0]               = IFP_oran_lphy_ctrl.ul_fft_scaler[0][3:0];
	assign IFP_oran_lphy_ctrl_new[0].ul_fft_scaler[1][3:0]               = IFP_oran_lphy_ctrl.ul_fft_scaler[1][3:0];	
    assign IFP_oran_lphy_ctrl_new[0].ul_fft_fraction_gain[0][15:0]       = IFP_oran_lphy_ctrl.ul_fft_fraction_gain[0][15:0];
	assign IFP_oran_lphy_ctrl_new[0].ul_fft_fraction_gain[1][15:0]       = IFP_oran_lphy_ctrl.ul_fft_fraction_gain[1][15:0];
    assign IFP_oran_lphy_ctrl_new[0].prach_en[0][3:0]                    = IFP_oran_lphy_ctrl.prach_en[0][3:0];
    assign IFP_oran_lphy_ctrl_new[0].prach_en[1][3:0]                    = IFP_oran_lphy_ctrl.prach_en[1][3:0];
    assign IFP_oran_lphy_ctrl_new[0].prach_format[0][3:0]                = IFP_oran_lphy_ctrl.prach_format[0][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_format[1][3:0]                = IFP_oran_lphy_ctrl.prach_format[1][3:0];
    assign IFP_oran_lphy_ctrl_new[0].prach_cp[0][15:0]                   = IFP_oran_lphy_ctrl.prach_cp[0][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_cp[1][15:0]                   = IFP_oran_lphy_ctrl.prach_cp[1][15:0];
    assign IFP_oran_lphy_ctrl_new[0].prach_use_sec_type3_freq_offset     = IFP_oran_lphy_ctrl.prach_use_sec_type3_freq_offset;
    assign IFP_oran_lphy_ctrl_new[0].prach_car_nco_lsb[0][31:0]          = IFP_oran_lphy_ctrl.prach_car_nco_lsb[0][31:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_car_nco_lsb[1][31:0]          = IFP_oran_lphy_ctrl.prach_car_nco_lsb[1][31:0];
    assign IFP_oran_lphy_ctrl_new[0].prach_car_nco_msb[0][6:0]           = IFP_oran_lphy_ctrl.prach_car_nco_msb[0][6:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_car_nco_msb[1][6:0]           = IFP_oran_lphy_ctrl.prach_car_nco_msb[1][6:0];
    assign IFP_oran_lphy_ctrl_new[0].prach_car_nco_sign[0]               = IFP_oran_lphy_ctrl.prach_car_nco_sign[0];
	assign IFP_oran_lphy_ctrl_new[0].prach_car_nco_sign[1]               = IFP_oran_lphy_ctrl.prach_car_nco_sign[1];	
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[0][0]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[0][1]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][1];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[0][2]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][2];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[0][3]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][3];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[1][0]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[1][1]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][1];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[1][2]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][2];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler_sign[1][3]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][3];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[0][0][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][0][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[0][1][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][1][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[0][2][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][2][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[0][3][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][3][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[1][0][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][0][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[1][1][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][1][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[1][2][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][2][3:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_scaler[1][3][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][3][3:0];	
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[0][0][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][0][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[0][1][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][1][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[0][2][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][2][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[0][3][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][3][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[1][0][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][0][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[1][1][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][1][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[1][2][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][2][15:0];
	assign IFP_oran_lphy_ctrl_new[0].prach_gain_fraction[1][3][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][3][15:0];		
    assign IFP_oran_lphy_ctrl_new[0].ul_lphy_oran_clear                  = IFP_oran_lphy_ctrl.ul_lphy_oran_clear;
    assign IFP_oran_lphy_ctrl_new[0].ul_lphy_oran_fifo_reset             = IFP_oran_lphy_ctrl.ul_lphy_oran_fifo_reset;
    assign IFP_oran_lphy_ctrl_new[0].prach_oran_clear                    = IFP_oran_lphy_ctrl.prach_oran_clear;
    assign IFP_oran_lphy_ctrl_new[0].prach_oran_fifo_reset               = IFP_oran_lphy_ctrl.prach_oran_fifo_reset;	
    assign IFP_oran_lphy_ctrl_new[0].lphy_oran_dbg_clear                 = IFP_oran_lphy_ctrl.lphy_oran_dbg_clear;
    assign IFP_oran_lphy_ctrl_new[0].lphy_oran_dbg_click                 = IFP_oran_lphy_ctrl.lphy_oran_dbg_click;
	
	
	assign IFP_oran_lphy_ctrl_new[1].dl_swap_ifft                        = IFP_oran_lphy_ctrl.dl_swap_ifft;
	assign IFP_oran_lphy_ctrl_new[1].ul_swap_fft                         = IFP_oran_lphy_ctrl.ul_swap_fft;	
	assign IFP_oran_lphy_ctrl_new[1].prach_swap_fft                      = IFP_oran_lphy_ctrl.prach_swap_fft;	
	assign IFP_oran_lphy_ctrl_new[1].dl_iq_endianness                    = IFP_oran_lphy_ctrl.dl_iq_endianness;
	assign IFP_oran_lphy_ctrl_new[1].ul_iq_endianness                    = IFP_oran_lphy_ctrl.ul_iq_endianness;	
	assign IFP_oran_lphy_ctrl_new[1].prach_iq_endianness                 = IFP_oran_lphy_ctrl.prach_iq_endianness;
    assign IFP_oran_lphy_ctrl_new[1].dl_ifft_gain_override[0]            = IFP_oran_lphy_ctrl.dl_ifft_gain_override[0];
    assign IFP_oran_lphy_ctrl_new[1].dl_ifft_gain_override[1]            = IFP_oran_lphy_ctrl.dl_ifft_gain_override[1];	
    assign IFP_oran_lphy_ctrl_new[1].ul_fft_gain_override[0]             = IFP_oran_lphy_ctrl.ul_fft_gain_override[0];
    assign IFP_oran_lphy_ctrl_new[1].ul_fft_gain_override[1]             = IFP_oran_lphy_ctrl.ul_fft_gain_override[1];	
	assign IFP_oran_lphy_ctrl_new[1].dl_route_c0_to_c1                   = IFP_oran_lphy_ctrl.dl_route_c0_to_c1;
    assign IFP_oran_lphy_ctrl_new[1].dl_lte_5g[0]                        = IFP_oran_lphy_ctrl.dl_lte_5g[0];
	assign IFP_oran_lphy_ctrl_new[1].dl_lte_5g[1]                        = IFP_oran_lphy_ctrl.dl_lte_5g[1];
    assign IFP_oran_lphy_ctrl_new[1].dl_extended_cp[0]                   = IFP_oran_lphy_ctrl.dl_extended_cp[0];
	assign IFP_oran_lphy_ctrl_new[1].dl_extended_cp[1]                   = IFP_oran_lphy_ctrl.dl_extended_cp[1];
    assign IFP_oran_lphy_ctrl_new[1].dl_cc_numerology[0][3:0]            = IFP_oran_lphy_ctrl.dl_cc_numerology[0][3:0];
	assign IFP_oran_lphy_ctrl_new[1].dl_cc_numerology[1][3:0]            = IFP_oran_lphy_ctrl.dl_cc_numerology[1][3:0];
    assign IFP_oran_lphy_ctrl_new[1].dl_ifft_scaler_sign[0]              = IFP_oran_lphy_ctrl.dl_ifft_scaler_sign[0];
	assign IFP_oran_lphy_ctrl_new[1].dl_ifft_scaler_sign[1]              = IFP_oran_lphy_ctrl.dl_ifft_scaler_sign[1];
    assign IFP_oran_lphy_ctrl_new[1].dl_ifft_scaler[0][3:0]              = IFP_oran_lphy_ctrl.dl_ifft_scaler[0][3:0];
	assign IFP_oran_lphy_ctrl_new[1].dl_ifft_scaler[1][3:0]              = IFP_oran_lphy_ctrl.dl_ifft_scaler[1][3:0];
    assign IFP_oran_lphy_ctrl_new[1].dl_ifft_fraction_gain[0][15:0]      = IFP_oran_lphy_ctrl.dl_ifft_fraction_gain[0][15:0];
	assign IFP_oran_lphy_ctrl_new[1].dl_ifft_fraction_gain[1][15:0]      = IFP_oran_lphy_ctrl.dl_ifft_fraction_gain[1][15:0];
    assign IFP_oran_lphy_ctrl_new[1].ul_lte_5g[0]                        = IFP_oran_lphy_ctrl.ul_lte_5g[0];
	assign IFP_oran_lphy_ctrl_new[1].ul_lte_5g[1]                        = IFP_oran_lphy_ctrl.ul_lte_5g[1];
    assign IFP_oran_lphy_ctrl_new[1].ul_extended_cp[0]                   = IFP_oran_lphy_ctrl.ul_extended_cp[0];
	assign IFP_oran_lphy_ctrl_new[1].ul_extended_cp[1]                   = IFP_oran_lphy_ctrl.ul_extended_cp[1];
    assign IFP_oran_lphy_ctrl_new[1].ul_cc_numerology[0][3:0]            = IFP_oran_lphy_ctrl.ul_cc_numerology[0][3:0];
	assign IFP_oran_lphy_ctrl_new[1].ul_cc_numerology[1][3:0]            = IFP_oran_lphy_ctrl.ul_cc_numerology[1][3:0];
    assign IFP_oran_lphy_ctrl_new[1].ul_fft_scaler_sign[0]               = IFP_oran_lphy_ctrl.ul_fft_scaler_sign[0];
	assign IFP_oran_lphy_ctrl_new[1].ul_fft_scaler_sign[1]               = IFP_oran_lphy_ctrl.ul_fft_scaler_sign[1];
    assign IFP_oran_lphy_ctrl_new[1].ul_fft_scaler[0][3:0]               = IFP_oran_lphy_ctrl.ul_fft_scaler[0][3:0];
	assign IFP_oran_lphy_ctrl_new[1].ul_fft_scaler[1][3:0]               = IFP_oran_lphy_ctrl.ul_fft_scaler[1][3:0];
    assign IFP_oran_lphy_ctrl_new[1].ul_fft_fraction_gain[0][15:0]       = IFP_oran_lphy_ctrl.ul_fft_fraction_gain[0][15:0];
	assign IFP_oran_lphy_ctrl_new[1].ul_fft_fraction_gain[1][15:0]       = IFP_oran_lphy_ctrl.ul_fft_fraction_gain[1][15:0];	
    assign IFP_oran_lphy_ctrl_new[1].prach_en[0][3:0]                    = IFP_oran_lphy_ctrl.prach_en[0][7:4];
    assign IFP_oran_lphy_ctrl_new[1].prach_en[1][3:0]                    = IFP_oran_lphy_ctrl.prach_en[1][7:4];
    assign IFP_oran_lphy_ctrl_new[1].prach_format[0][3:0]                = IFP_oran_lphy_ctrl.prach_format[0][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_format[1][3:0]                = IFP_oran_lphy_ctrl.prach_format[1][3:0];
    assign IFP_oran_lphy_ctrl_new[1].prach_cp[0][15:0]                   = IFP_oran_lphy_ctrl.prach_cp[0][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_cp[1][15:0]                   = IFP_oran_lphy_ctrl.prach_cp[1][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_use_sec_type3_freq_offset     = IFP_oran_lphy_ctrl.prach_use_sec_type3_freq_offset;
    assign IFP_oran_lphy_ctrl_new[1].prach_car_nco_lsb[0][31:0]          = IFP_oran_lphy_ctrl.prach_car_nco_lsb[0][31:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_car_nco_lsb[1][31:0]          = IFP_oran_lphy_ctrl.prach_car_nco_lsb[1][31:0];
    assign IFP_oran_lphy_ctrl_new[1].prach_car_nco_msb[0][6:0]           = IFP_oran_lphy_ctrl.prach_car_nco_msb[0][6:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_car_nco_msb[1][6:0]           = IFP_oran_lphy_ctrl.prach_car_nco_msb[1][6:0];
    assign IFP_oran_lphy_ctrl_new[1].prach_car_nco_sign[0]               = IFP_oran_lphy_ctrl.prach_car_nco_sign[0];
	assign IFP_oran_lphy_ctrl_new[1].prach_car_nco_sign[1]               = IFP_oran_lphy_ctrl.prach_car_nco_sign[1];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[0][0]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[0][1]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][1];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[0][2]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][2];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[0][3]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[0][3];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[1][0]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[1][1]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][1];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[1][2]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][2];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler_sign[1][3]        = IFP_oran_lphy_ctrl.prach_gain_scaler_sign[1][3];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[0][0][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][4][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[0][1][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][5][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[0][2][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][6][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[0][3][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[0][7][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[1][0][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][4][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[1][1][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][5][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[1][2][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][6][3:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_scaler[1][3][3:0]        = IFP_oran_lphy_ctrl.prach_gain_scaler[1][7][3:0];	
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[0][0][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][4][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[0][1][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][5][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[0][2][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][6][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[0][3][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[0][7][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[1][0][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][4][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[1][1][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][5][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[1][2][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][6][15:0];
	assign IFP_oran_lphy_ctrl_new[1].prach_gain_fraction[1][3][15:0]     = IFP_oran_lphy_ctrl.prach_gain_fraction[1][7][15:0];	
	assign IFP_oran_lphy_ctrl_new[1].ul_lphy_oran_clear                  = IFP_oran_lphy_ctrl.ul_lphy_oran_clear;
	assign IFP_oran_lphy_ctrl_new[1].ul_lphy_oran_fifo_reset             = IFP_oran_lphy_ctrl.ul_lphy_oran_fifo_reset;	
	assign IFP_oran_lphy_ctrl_new[1].prach_oran_clear                    = IFP_oran_lphy_ctrl.prach_oran_clear;
	assign IFP_oran_lphy_ctrl_new[1].prach_oran_fifo_reset               = IFP_oran_lphy_ctrl.prach_oran_fifo_reset;
	assign IFP_oran_lphy_ctrl_new[1].lphy_oran_dbg_clear                 = IFP_oran_lphy_ctrl.lphy_oran_dbg_clear;
	assign IFP_oran_lphy_ctrl_new[1].lphy_oran_dbg_click                 = IFP_oran_lphy_ctrl.lphy_oran_dbg_click;	
	
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_int_frac_delay_trig             = IFP_ul_dfe_ctrl.ul_ant_int_frac_delay_trig;
	assign IFP_ul_dfe_ctrl_new[0].ul_car_nco_lsb[0][31:0]                = IFP_ul_dfe_ctrl.ul_car_nco_lsb[0][31:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_car_nco_lsb[1][31:0]                = IFP_ul_dfe_ctrl.ul_car_nco_lsb[1][31:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_car_nco_msb[0][6:0]                 = IFP_ul_dfe_ctrl.ul_car_nco_msb[0][6:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_car_nco_msb[1][6:0]                 = IFP_ul_dfe_ctrl.ul_car_nco_msb[1][6:0];			
	assign IFP_ul_dfe_ctrl_new[0].ul_car_nco_msb[0][7]                   = IFP_ul_dfe_ctrl.ul_car_nco_sign[0];		
	assign IFP_ul_dfe_ctrl_new[0].ul_car_nco_msb[1][7]                   = IFP_ul_dfe_ctrl.ul_car_nco_sign[1];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler_sign[0][3:0]     = IFP_ul_dfe_ctrl.ul_stream_gain_scaler_sign[0][3:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler_sign[1][3:0]     = IFP_ul_dfe_ctrl.ul_stream_gain_scaler_sign[1][3:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[0][0][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][0][3:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[0][1][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][1][3:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[0][2][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][2][3:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[0][3][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][3][3:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[1][0][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][0][3:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[1][1][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][1][3:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[1][2][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][2][3:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_scaler[1][3][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][3][3:0];																	     
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[0][0][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][0][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[0][1][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][1][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[0][2][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][2][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[0][3][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][3][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[1][0][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][0][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[1][1][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][1][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[1][2][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][2][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_stream_gain_fraction[1][3][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][3][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_scaler_sign[3:0]           = IFP_ul_dfe_ctrl.ul_ant_gain_scaler_sign[3:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_scaler[0][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[0][3:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_scaler[1][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[1][3:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_scaler[2][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[2][3:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_scaler[3][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[3][3:0];		
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_fraction[0][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[0][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_fraction[1][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[1][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_fraction[2][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[2][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_ant_gain_fraction[3][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[3][15:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[0][0][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][0][6:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[0][1][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][1][6:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[0][2][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][2][6:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[0][3][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][3][6:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[1][0][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][0][6:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[1][1][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][1][6:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[1][2][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][2][6:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_int_delay[1][3][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][3][6:0];		
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[0][0][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][0][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[0][1][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][1][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[0][2][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][2][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[0][3][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][3][15:0];	
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[1][0][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][0][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[1][1][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][1][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[1][2][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][2][15:0];
	assign IFP_ul_dfe_ctrl_new[0].ul_frac_delay[1][3][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][3][15:0];	

	assign IFP_ul_dfe_ctrl_new[1].ul_ant_int_frac_delay_trig             = IFP_ul_dfe_ctrl.ul_ant_int_frac_delay_trig;
	assign IFP_ul_dfe_ctrl_new[1].ul_car_nco_lsb[0][31:0]                = IFP_ul_dfe_ctrl.ul_car_nco_lsb[0][31:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_car_nco_lsb[1][31:0]                = IFP_ul_dfe_ctrl.ul_car_nco_lsb[1][31:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_car_nco_msb[0][6:0]                 = IFP_ul_dfe_ctrl.ul_car_nco_msb[0][6:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_car_nco_msb[1][6:0]                 = IFP_ul_dfe_ctrl.ul_car_nco_msb[1][6:0];			
	assign IFP_ul_dfe_ctrl_new[1].ul_car_nco_msb[0][7]                   = IFP_ul_dfe_ctrl.ul_car_nco_sign[0];		
	assign IFP_ul_dfe_ctrl_new[1].ul_car_nco_msb[1][7]                   = IFP_ul_dfe_ctrl.ul_car_nco_sign[1];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler_sign[0][3:0]     = IFP_ul_dfe_ctrl.ul_stream_gain_scaler_sign[0][7:4];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler_sign[1][3:0]     = IFP_ul_dfe_ctrl.ul_stream_gain_scaler_sign[1][7:4];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[0][0][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][4][3:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[0][1][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][5][3:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[0][2][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][6][3:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[0][3][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[0][7][3:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[1][0][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][4][3:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[1][1][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][5][3:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[1][2][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][6][3:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_scaler[1][3][3:0]       = IFP_ul_dfe_ctrl.ul_stream_gain_scaler[1][7][3:0];																	     
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[0][0][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][4][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[0][1][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][5][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[0][2][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][6][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[0][3][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[0][7][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[1][0][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][4][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[1][1][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][5][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[1][2][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][6][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_stream_gain_fraction[1][3][15:0]    = IFP_ul_dfe_ctrl.ul_stream_gain_fraction[1][7][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_scaler_sign[3:0]           = IFP_ul_dfe_ctrl.ul_ant_gain_scaler_sign[7:4];	
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_scaler[0][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[4][3:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_scaler[1][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[5][3:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_scaler[2][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[6][3:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_scaler[3][3:0]             = IFP_ul_dfe_ctrl.ul_ant_gain_scaler[7][3:0];		
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_fraction[0][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[4][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_fraction[1][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[5][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_fraction[2][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[6][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_ant_gain_fraction[3][15:0]          = IFP_ul_dfe_ctrl.ul_ant_gain_fraction[7][15:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[0][0][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][4][6:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[0][1][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][5][6:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[0][2][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][6][6:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[0][3][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[0][7][6:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[1][0][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][4][6:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[1][1][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][5][6:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[1][2][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][6][6:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_int_delay[1][3][6:0]                = IFP_ul_dfe_ctrl.ul_int_delay[1][7][6:0];		
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[0][0][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][4][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[0][1][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][5][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[0][2][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][6][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[0][3][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[0][7][15:0];	
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[1][0][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][4][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[1][1][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][5][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[1][2][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][6][15:0];
	assign IFP_ul_dfe_ctrl_new[1].ul_frac_delay[1][3][15:0]              = IFP_ul_dfe_ctrl.ul_frac_delay[1][7][15:0];	
	
	logic  [7:0] s_dpd_tuser_field;	
	assign IFP_dpd_s_axis_din_new.tdata    = {IFP_dpd_s_axis_din[1].tdata, IFP_dpd_s_axis_din[0].tdata};
	assign IFP_dpd_s_axis_din_new.tlast    = IFP_dpd_s_axis_din[0].tlast | IFP_dpd_s_axis_din[1].tlast;
	assign IFP_dpd_s_axis_din[0].tready    = IFP_dpd_s_axis_din_new.tready;
	assign IFP_dpd_s_axis_din[1].tready    = IFP_dpd_s_axis_din_new.tready;
//	assign IFP_dpd_s_axis_din_new.tuser    = {IFP_dpd_s_axis_din[1].tuser,IFP_dpd_s_axis_din[0].tuser};
    assign s_dpd_tuser_field               = {4'd0,syn_data_dl_ul_5ms,syn_data_dl_ul_5ms,tuser_dl_frm_mrkr_10ms,1'b0};
	assign IFP_dpd_s_axis_din_new.tuser    = {8{s_dpd_tuser_field}};
	assign IFP_dpd_s_axis_din_new.tvalid   = IFP_dpd_s_axis_din[0].tvalid | IFP_dpd_s_axis_din[1].tvalid;
										   
	assign IFP_dpd_m_axis_dout_new.tready  = IFP_dpd_m_axis_dout[0].tready | IFP_dpd_m_axis_dout[1].tready;
	assign IFP_dpd_m_axis_dout[0].tdata    = IFP_dpd_m_axis_dout_new.tdata[127:0];
	assign IFP_dpd_m_axis_dout[0].tlast    = IFP_dpd_m_axis_dout_new.tlast;
	assign IFP_dpd_m_axis_dout[0].tuser    = IFP_dpd_m_axis_dout_new.tuser[31:0];
	assign IFP_dpd_m_axis_dout[0].tvalid   = IFP_dpd_m_axis_dout_new.tvalid;

	assign IFP_dpd_m_axis_dout[1].tdata    = IFP_dpd_m_axis_dout_new.tdata[255:128];
	assign IFP_dpd_m_axis_dout[1].tlast    = IFP_dpd_m_axis_dout_new.tlast;
	assign IFP_dpd_m_axis_dout[1].tuser    = IFP_dpd_m_axis_dout_new.tuser[63:32];
	assign IFP_dpd_m_axis_dout[1].tvalid   = IFP_dpd_m_axis_dout_new.tvalid;
										   
										   
	assign IFP_cfr_s_axis_din_new.tdata    = {IFP_cfr_s_axis_din[1].tdata, IFP_cfr_s_axis_din[0].tdata};
	assign IFP_cfr_s_axis_din_new.tlast    = IFP_cfr_s_axis_din[0].tlast | IFP_cfr_s_axis_din[1].tlast;
	assign IFP_cfr_s_axis_din[0].tready    = IFP_cfr_s_axis_din_new.tready;
	assign IFP_cfr_s_axis_din[1].tready    = IFP_cfr_s_axis_din_new.tready;
	assign IFP_cfr_s_axis_din_new.tuser    = IFP_cfr_s_axis_din[0].tuser;
	assign IFP_cfr_s_axis_din_new.tvalid   = IFP_cfr_s_axis_din[0].tvalid | IFP_cfr_s_axis_din[1].tvalid;	
	
	assign IFP_cfr_m_axis_dout_new.tready  = IFP_cfr_m_axis_dout[0].tready | IFP_cfr_m_axis_dout[1].tready;
	assign IFP_cfr_m_axis_dout[0].tdata    = IFP_cfr_m_axis_dout_new.tdata[127:0];
	assign IFP_cfr_m_axis_dout[0].tlast    = IFP_cfr_m_axis_dout_new.tlast;
	assign IFP_cfr_m_axis_dout[0].tuser    = IFP_cfr_m_axis_dout_new.tuser;
	assign IFP_cfr_m_axis_dout[0].tvalid   = IFP_cfr_m_axis_dout_new.tvalid;

	assign IFP_cfr_m_axis_dout[1].tdata    = IFP_cfr_m_axis_dout_new.tdata[255:128];
	assign IFP_cfr_m_axis_dout[1].tlast    = IFP_cfr_m_axis_dout_new.tlast;
	assign IFP_cfr_m_axis_dout[1].tuser    = IFP_cfr_m_axis_dout_new.tuser;
	assign IFP_cfr_m_axis_dout[1].tvalid   = IFP_cfr_m_axis_dout_new.tvalid;	
	
	
	
	
	
endmodule
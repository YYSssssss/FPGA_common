

module jb_dl_dfe_input_waveform #(
   parameter PTR_WIDTH =15,
   parameter PRECISION =16
) (
   input 				clk_en,
   input 				clk,
   input 				resetn,
   input 				IFP_iwavebuf_porta_rst,
   input 				IFP_iwavebuf_porta_clk, 
					jb_ram_sp_if.mem IFP_iwavebuf_porta,

   input [PTR_WIDTH-1:0] 		ptr,
   input [2*PRECISION-1:0] 		dina,
   input [3:0]                          wea,


   output logic signed [PRECISION-1 :0] real_value,
   output logic signed [PRECISION-1 :0] imag_value

 );

   logic [2*PRECISION-1:0] 	  douta;
   logic [PTR_WIDTH-1:0] 		ptr_reg;
   logic [2*PRECISION-1:0] 	  dina_reg;
   logic [2*PRECISION-1:0] 	  wea_reg;
   
   
     always @(posedge clk) begin
      if (!resetn) begin
	 ptr_reg<= 0;
	 wea_reg <= 0;
	 dina_reg <=0;
      end
      else if (clk_en) begin
	 ptr_reg<= ptr;
	 wea_reg <= wea;
	 dina_reg <=dina;
	 
      end
    end // always @ (posedge clk)

/*
      logic bram_porta_en;
      assign bram_porta_en = clk_en;
*/

// bram_iwaveform bram_input_waveform (
//  .clka(clk),    // input wire clka
//  //.ena (bram_porta_en),
//  .wea(wea_reg),
//  .addra({{(32-PTR_WIDTH){1'b0}},ptr_reg,2'b00}),  // input wire [31 : 0] addra
//  .dina(dina_reg),
//  .douta(douta),  // output wire [31 : 0] douta
//  .clkb(IFP_iwavebuf_porta_clk),
//  .rstb(IFP_iwavebuf_porta_rst),
//  .enb(IFP_iwavebuf_porta.en),
//  .web(IFP_iwavebuf_porta.wr_en),
//  .addrb(IFP_iwavebuf_porta.addr),     // input wire [14:0] addr
//  .dinb(IFP_iwavebuf_porta.wr_data),   // input wire [31:0] din
//  .doutb(IFP_iwavebuf_porta.rd_data)   // input wire [31:0] dout
//);

   /*
  always @(posedge clk) begin
       real_value<=  $signed(douta[PRECISION-1:0]);
       imag_value<=  $signed(douta[2*PRECISION-1:PRECISION]);
    end // always @ (posedge clk)
*/
   

      assign real_value =  $signed(douta[PRECISION-1:0]);
      assign imag_value =  $signed(douta[2*PRECISION-1:PRECISION]);
/*
always @(*) begin
   real_value= 0;
   imag_value=0;
    case(ptr)
    0    : begin
              real_value= 0;
              imag_value=0;
            end
    1     : begin
              real_value= 0;
              imag_value=0;
            end
    2     : begin
              real_value= 0;
              imag_value=0;
            end
    3     : begin
              real_value= 0;
              imag_value=0;
            end
    4     : begin
              real_value= 0;
              imag_value=0;
            end
    5     : begin
              real_value= 0;
              imag_value=0;
            end
    6     : begin
              real_value= 0;
              imag_value=0;
            end
    7     : begin
              real_value= 0;
              imag_value=0;
            end
    8     : begin
              real_value= 0;
              imag_value=0;
            end
    9     : begin
              real_value= 0;
              imag_value=0;
            end
    10     : begin
              real_value= 0;
              imag_value=0;
            end
    11    : begin
              real_value= 0;
              imag_value=0;
            end
    12    : begin
              real_value= 0;
              imag_value=0;
            end
    13    : begin
              real_value= 0;
              imag_value=0;
            end
    14    : begin
              real_value= 0;
              imag_value=0;
            end
    15    : begin
              real_value= 1;
              imag_value=0;
            end
    16    : begin
              real_value= -2;
              imag_value=0;
            end
    17    : begin
              real_value= 0;
              imag_value=0;
            end
    18    : begin
              real_value= 3;
              imag_value=0;
            end
    19    : begin
              real_value= -3;
              imag_value=0;
            end
    20    : begin
              real_value= -3;
              imag_value=0;
            end
    21    : begin
              real_value= 7;
              imag_value=0;
            end
    22    : begin
              real_value= 0;
              imag_value=0;
            end
    23    : begin
              real_value= -9;
              imag_value=0;
            end
    24    : begin
              real_value= 8;
              imag_value=0;
            end
    25    : begin
              real_value= 6;
              imag_value=0;
            end
    26    : begin
              real_value= -15;
              imag_value=1;
            end
    27    : begin
              real_value= 3;
              imag_value=0;
            end
    28    : begin
              real_value= 16;
              imag_value=0;
            end
    29    : begin
              real_value= -18;
              imag_value=2;
            end
    30    : begin
              real_value= -6;
              imag_value=0;
            end
    31    : begin
              real_value= 28;
              imag_value=-1;
            end
    32    : begin
              real_value= -12;
              imag_value=3;
            end
    33    : begin
              real_value= -25;
              imag_value=0;
            end
    34    : begin
              real_value= 36;
              imag_value=-3;
            end
    35    : begin
              real_value= 4;
              imag_value=2;
            end
    36    : begin
              real_value= -46;
              imag_value=3;
            end
    37    : begin
              real_value= 30;
              imag_value=-4;
            end
    38    : begin
              real_value= 33;
              imag_value=0;
            end
    39    : begin
              real_value= -63;
              imag_value=7;
            end
    40    : begin
              real_value= 4;
              imag_value=-3;
            end
    41    : begin
              real_value= 71;
              imag_value=-2;
            end
    42    : begin
              real_value= -60;
              imag_value=10;
            end
    43    : begin
              real_value= -40;
              imag_value=0;
            end
    44    : begin
              real_value= 101;
              imag_value=-8;
            end
    45    : begin
              real_value= -28;
              imag_value=10;
            end
    46    : begin
              real_value= -100;
              imag_value=4;
            end
    47    : begin
              real_value= 107;
              imag_value=-14;
            end
    48    : begin
              real_value= 36;
              imag_value=5;
            end
    49    : begin
              real_value= -156;
              imag_value=12;
            end
    50    : begin
              real_value= 70;
              imag_value=-17;
            end
    51    : begin
              real_value= 129;
              imag_value=-2;
            end
    52    : begin
              real_value= -183;
              imag_value=22;
            end
    53    : begin
              real_value= -18;
              imag_value=-13;
            end
    54    : begin
              real_value= 229;
              imag_value=-17;
            end
    55    : begin
              real_value= -149;
              imag_value=27;
            end
    56    : begin
              real_value= -159;
              imag_value=-1;
            end
    57    : begin
              real_value= 299;
              imag_value=-33;
            end
    58    : begin
              real_value= -30;
              imag_value=25;
            end
    59    : begin
              real_value= -331;
              imag_value=18;
            end
    60    : begin
              real_value= 292;
              imag_value=-47;
            end
    61    : begin
              real_value= 183;
              imag_value=11;
            end
    62    : begin
              real_value= -493;
              imag_value=48;
            end
    63    : begin
              real_value= 156;
              imag_value=-50;
            end
    64    : begin
              real_value= 501;
              imag_value=-17;
            end
    65    : begin
              real_value= -587;
              imag_value=82;
            end
    66    : begin
              real_value= -178;
              imag_value=-36;
            end
    67    : begin
              real_value= 933;
              imag_value=-72;
            end
    68    : begin
              real_value= -525;
              imag_value=117;
            end
    69    : begin
              real_value= -902;
              imag_value=7;
            end
    70    : begin
              real_value= 1648;
              imag_value=-174;
            end
    71    : begin
              real_value= -65;
              imag_value=162;
            end
    72    : begin
              real_value= -3446;
              imag_value=145;
            end
    73    : begin
              real_value= 6382;
              imag_value=-555;
            end
    74    : begin
              real_value= 26397;
              imag_value=750;
            end
    75    : begin
              real_value= 32766;
              imag_value=6097;
            end
    76    : begin
              real_value= 30155;
              imag_value=13177;
            end
    77    : begin
              real_value= 25133;
              imag_value=19027;
            end
    78    : begin
              real_value= 23281;
              imag_value=23736;
            end
    79    : begin
              real_value= 17611;
              imag_value=27970;
            end
    80    : begin
              real_value= 10106;
              imag_value=30964;
            end
    81    : begin
              real_value= 4708;
              imag_value=32371;
            end
    82    : begin
              real_value= -1549;
              imag_value=32653;
            end
    83    : begin
              real_value= -9232;
              imag_value=31659;
            end
    84    : begin
              real_value= -15133;
              imag_value=29123;
            end
    85    : begin
              real_value= -20081;
              imag_value=25442;
            end
    86    : begin
              real_value= -25503;
              imag_value=20833;
            end
    87    : begin
              real_value= -29314;
              imag_value=15218;
            end
    88    : begin
              real_value= -31172;
              imag_value=8947;
            end
    89    : begin
              real_value= -32636;
              imag_value=2428;
            end
    90    : begin
              real_value= -32767;
              imag_value=-4249;
            end
    91    : begin
              real_value= -30778;
              imag_value=-10818;
            end
    92    : begin
              real_value= -27946;
              imag_value=-16844;
            end
    93    : begin
              real_value= -24322;
              imag_value=-22170;
            end
    94    : begin
              real_value= -19065;
              imag_value=-26648;
            end
    95    : begin
              real_value= -13089;
              imag_value=-29965;
            end
    96    : begin
              real_value= -7044;
              imag_value=-31999;
            end
    97    : begin
              real_value= -341;
              imag_value=-32763;
            end
    98    : begin
              real_value= 6547;
              imag_value=-32149;
            end
    99    : begin
              real_value= 12749;
              imag_value=-30149;
            end
    100    : begin
              real_value= 18535;
              imag_value=-26931;
            end
    101   : begin
              real_value= 23827;
              imag_value=-22605;
            end
    102   : begin
              real_value= 27851;
              imag_value=-17294;
            end
    103   : begin
              real_value= 30652;
              imag_value=-11277;
            end
    104   : begin
              real_value= 32447;
              imag_value=-4816;
            end
    105   : begin
              real_value= 32766;
              imag_value=1873;
            end
    106   : begin
              real_value= 31573;
              imag_value=8488;
            end
    107   : begin
              real_value= 29257;
              imag_value=14724;
            end
    108   : begin
              real_value= 25725;
              imag_value=20360;
            end
    109   : begin
              real_value= 20954;
              imag_value=25162;
            end
    110   : begin
              real_value= 15411;
              imag_value=28893;
            end
    111   : begin
              real_value= 9300;
              imag_value=31421;
            end
    112   : begin
              real_value= 2671;
              imag_value=32656;
            end
    113   : begin
              real_value= -4046;
              imag_value=32518;
            end
    114   : begin
              real_value= -10504;
              imag_value=31018;
            end
    115   : begin
              real_value= -16597;
              imag_value=28238;
            end
    116   : begin
              real_value= -22030;
              imag_value=24278;
            end
    117   : begin
              real_value= -26465;
              imag_value=19297;
            end
    118   : begin
              real_value= -29821;
              imag_value=13520;
            end
    119   : begin
              real_value= -31983;
              imag_value=7181;
            end
    120   : begin
              real_value= -32762;
              imag_value=534;
            end
    121   : begin
              real_value= -32167;
              imag_value=-6128;
            end
    122   : begin
              real_value= -30274;
              imag_value=-12535;
            end
    123   : begin
              real_value= -27099;
              imag_value=-18422;
            end
    124   : begin
              real_value= -22772;
              imag_value=-23542;
            end
    125   : begin
              real_value= -17525;
              imag_value=-27677;
            end
    126   : begin
              real_value= -11547;
              imag_value=-30660;
            end
    127   : begin
              real_value= -5067;
              imag_value=-32366;
            end
    128   : begin
              real_value= 1610;
              imag_value=-32720;
            end
    129   : begin
              real_value= 8214;
              imag_value=-31711;
            end
    130   : begin
              real_value= 14490;
              imag_value=-29381;
            end
    131   : begin
              real_value= 20158;
              imag_value=-25826;
            end
    132   : begin
              real_value= 24978;
              imag_value=-21193;
            end
    133   : begin
              real_value= 28764;
              imag_value=-15678;
            end
    134   : begin
              real_value= 31352;
              imag_value=-9508;
            end
    135   : begin
              real_value= 32627;
              imag_value=-2942;
            end
    136   : begin
              real_value= 32545;
              imag_value=3743;
            end
    137   : begin
              real_value= 31108;
              imag_value=10275;
            end
    138   : begin
              real_value= 28371;
              imag_value=16380;
            end
    139   : begin
              real_value= 24452;
              imag_value=21801;
            end
    140   : begin
              real_value= 19515;
              imag_value=26314;
            end
    141   : begin
              real_value= 13764;
              imag_value=29729;
            end
    142   : begin
              real_value= 7438;
              imag_value=31905;
            end
    143   : begin
              real_value= 802;
              imag_value=32750;
            end
    144   : begin
              real_value= -5864;
              imag_value=32231;
            end
    145   : begin
              real_value= -12288;
              imag_value=30369;
            end
    146   : begin
              real_value= -18200;
              imag_value=27240;
            end
    147   : begin
              real_value= -23354;
              imag_value=22974;
            end
    148   : begin
              real_value= -27534;
              imag_value=17752;
            end
    149   : begin
              real_value= -30565;
              imag_value=11790;
            end
    150   : begin
              real_value= -32323;
              imag_value=5336;
            end
    151   : begin
              real_value= -32733;
              imag_value=-1338;
            end
    152   : begin
              real_value= -31779;
              imag_value=-7959;
            end
    153   : begin
              real_value= -29499;
              imag_value=-14248;
            end
    154   : begin
              real_value= -25990;
              imag_value=-19943;
            end
    155   : begin
              real_value= -21399;
              imag_value=-24806;
            end
    156   : begin
              real_value= -15914;
              imag_value=-28636;
            end
    157   : begin
              real_value= -9765;
              imag_value=-31271;
            end
    158   : begin
              real_value= -3210;
              imag_value=-32603;
            end
    159   : begin
              real_value= 3476;
              imag_value=-32575;
            end
    160   : begin
              real_value= 10021;
              imag_value=-31191;
            end
    161   : begin
              real_value= 16148;
              imag_value=-28506;
            end
    162   : begin
              real_value= 21600;
              imag_value=-24630;
            end
    163   : begin
              real_value= 26152;
              imag_value=-19729;
            end
    164   : begin
              real_value= 29615;
              imag_value=-14006;
            end
    165   : begin
              real_value= 31843;
              imag_value=-7699;
            end
    166   : begin
              real_value= 32743;
              imag_value=-1070;
            end
    167   : begin
              real_value= 32278;
              imag_value=5599;
            end
    168   : begin
              real_value= 30468;
              imag_value=12039;
            end
    169   : begin
              real_value= 27387;
              imag_value=17977;
            end
    170   : begin
              real_value= 23165;
              imag_value=23165;
            end
    171   : begin
              real_value= 17977;
              imag_value=27387;
            end
    172   : begin
              real_value= 12039;
              imag_value=30468;
            end
    173   : begin
              real_value= 5599;
              imag_value=32278;
            end
    174   : begin
              real_value= -1070;
              imag_value=32743;
            end
    175   : begin
              real_value= -7699;
              imag_value=31843;
            end
    176   : begin
              real_value= -14006;
              imag_value=29615;
            end
    177   : begin
              real_value= -19729;
              imag_value=26152;
            end
    178   : begin
              real_value= -24630;
              imag_value=21600;
            end
    179   : begin
              real_value= -28506;
              imag_value=16148;
            end
    180   : begin
              real_value= -31191;
              imag_value=10021;
            end
    181   : begin
              real_value= -32575;
              imag_value=3476;
            end
    182   : begin
              real_value= -32603;
              imag_value=-3210;
            end
    183   : begin
              real_value= -31271;
              imag_value=-9765;
            end
    184   : begin
              real_value= -28636;
              imag_value=-15914;
            end
    185   : begin
              real_value= -24806;
              imag_value=-21399;
            end
    186   : begin
              real_value= -19943;
              imag_value=-25990;
            end
    187   : begin
              real_value= -14248;
              imag_value=-29499;
            end
    188   : begin
              real_value= -7959;
              imag_value=-31779;
            end
    189   : begin
              real_value= -1338;
              imag_value=-32733;
            end
    190   : begin
              real_value= 5336;
              imag_value=-32323;
            end
    191   : begin
              real_value= 11790;
              imag_value=-30565;
            end
    192   : begin
              real_value= 17752;
              imag_value=-27534;
            end
    193   : begin
              real_value= 22974;
              imag_value=-23354;
            end
    194   : begin
              real_value= 27240;
              imag_value=-18200;
            end
    195   : begin
              real_value= 30369;
              imag_value=-12288;
            end
    196   : begin
              real_value= 32231;
              imag_value=-5864;
            end
    197   : begin
              real_value= 32750;
              imag_value=802;
            end
    198   : begin
              real_value= 31905;
              imag_value=7438;
            end
    199   : begin
              real_value= 29729;
              imag_value=13764;
            end
    200   : begin
              real_value= 26314;
              imag_value=19515;
            end
    201   : begin
              real_value= 21801;
              imag_value=24453;
            end
    202   : begin
              real_value= 16380;
              imag_value=28371;
            end
    203   : begin
              real_value= 10275;
              imag_value=31107;
            end
    204   : begin
              real_value= 3742;
              imag_value=32547;
            end
    205   : begin
              real_value= -2942;
              imag_value=32629;
            end
    206   : begin
              real_value= -9508;
              imag_value=31351;
            end
    207   : begin
              real_value= -15678;
              imag_value=28766;
            end
    208   : begin
              real_value= -21194;
              imag_value=24981;
            end
    209   : begin
              real_value= -25826;
              imag_value=20154;
            end
    210   : begin
              real_value= -29382;
              imag_value=14489;
            end
    211   : begin
              real_value= -31713;
              imag_value=8219;
            end
    212   : begin
              real_value= -32721;
              imag_value=1606;
            end
    213   : begin
              real_value= -32365;
              imag_value=-5071;
            end
    214   : begin
              real_value= -30661;
              imag_value=-11539;
            end
    215   : begin
              real_value= -27678;
              imag_value=-17525;
            end
    216   : begin
              real_value= -23541;
              imag_value=-22782;
            end
    217   : begin
              real_value= -18423;
              imag_value=-27090;
            end
    218   : begin
              real_value= -12537;
              imag_value=-30267;
            end
    219   : begin
              real_value= -6127;
              imag_value=-32183;
            end
    220   : begin
              real_value= 535;
              imag_value=-32757;
            end
    221   : begin
              real_value= 7177;
              imag_value=-31965;
            end
    222   : begin
              real_value= 13520;
              imag_value=-29841;
            end
    223   : begin
              real_value= 19299;
              imag_value=-26472;
            end
    224   : begin
              real_value= 24274;
              imag_value=-22001;
            end
    225   : begin
              real_value= 28236;
              imag_value=-16611;
            end
    226   : begin
              real_value= 31023;
              imag_value=-10529;
            end
    227   : begin
              real_value= 32515;
              imag_value=-4009;
            end
    228   : begin
              real_value= 32651;
              imag_value=2676;
            end
    229   : begin
              real_value= 31426;
              imag_value=9253;
            end
    230   : begin
              real_value= 28892;
              imag_value=15442;
            end
    231   : begin
              real_value= 25154;
              imag_value=20988;
            end
    232   : begin
              real_value= 20365;
              imag_value=25661;
            end
    233   : begin
              real_value= 14728;
              imag_value=29263;
            end
    234   : begin
              real_value= 8477;
              imag_value=31645;
            end
    235   : begin
              real_value= 1874;
              imag_value=32707;
            end
    236   : begin
              real_value= -4806;
              imag_value=32407;
            end
    237   : begin
              real_value= -11289;
              imag_value=30755;
            end
    238   : begin
              real_value= -17299;
              imag_value=27820;
            end
    239   : begin
              real_value= -22589;
              imag_value=23726;
            end
    240   : begin
              real_value= -26938;
              imag_value=18644;
            end
    241   : begin
              real_value= -30163;
              imag_value=12784;
            end
    242   : begin
              real_value= -32131;
              imag_value=6390;
            end
    243   : begin
              real_value= -32759;
              imag_value=-267;
            end
    244   : begin
              real_value= -32022;
              imag_value=-6915;
            end
    245   : begin
              real_value= -29950;
              imag_value=-13274;
            end
    246   : begin
              real_value= -26630;
              imag_value=-19081;
            end
    247   : begin
              real_value= -22199;
              imag_value=-24092;
            end
    248   : begin
              real_value= -16842;
              imag_value=-28100;
            end
    249   : begin
              real_value= -10783;
              imag_value=-30935;
            end
    250   : begin
              real_value= -4275;
              imag_value=-32481;
            end
    251   : begin
              real_value= 2408;
              imag_value=-32673;
            end
    252   : begin
              real_value= 8995;
              imag_value=-31501;
            end
    253   : begin
              real_value= 15206;
              imag_value=-29017;
            end
    254   : begin
              real_value= 20783;
              imag_value=-25324;
            end
    255   : begin
              real_value= 25494;
              imag_value=-20575;
            end
    256   : begin
              real_value= 29142;
              imag_value=-14968;
            end
    257   : begin
              real_value= 31575;
              imag_value=-8737;
            end
    258   : begin
              real_value= 32691;
              imag_value=-2142;
            end
    259   : begin
              real_value= 32445;
              imag_value=4540;
            end
    260   : begin
              real_value= 30846;
              imag_value=11036;
            end
    261   : begin
              real_value= 27961;
              imag_value=17072;
            end
    262   : begin
              real_value= 23911;
              imag_value=22395;
            end
    263   : begin
              real_value= 18863;
              imag_value=26784;
            end
    264   : begin
              real_value= 13030;
              imag_value=30057;
            end
    265   : begin
              real_value= 6654;
              imag_value=32077;
            end
    266   : begin
              real_value= 0;
              imag_value=32760;
            end
    267   : begin
              real_value= -6654;
              imag_value=32077;
            end
    268   : begin
              real_value= -13030;
              imag_value=30057;
            end
    269   : begin
              real_value= -18863;
              imag_value=26784;
            end
    270   : begin
              real_value= -23911;
              imag_value=22395;
            end
    271   : begin
              real_value= -27961;
              imag_value=17072;
            end
    272   : begin
              real_value= -30846;
              imag_value=11036;
            end
    273   : begin
              real_value= -32445;
              imag_value=4540;
            end
    274   : begin
              real_value= -32691;
              imag_value=-2142;
            end
    275   : begin
              real_value= -31575;
              imag_value=-8737;
            end
    276   : begin
              real_value= -29142;
              imag_value=-14968;
            end
    277   : begin
              real_value= -25494;
              imag_value=-20575;
            end
    278   : begin
              real_value= -20783;
              imag_value=-25324;
            end
    279   : begin
              real_value= -15206;
              imag_value=-29017;
            end
    280   : begin
              real_value= -8995;
              imag_value=-31501;
            end
    281   : begin
              real_value= -2408;
              imag_value=-32673;
            end
    282   : begin
              real_value= 4275;
              imag_value=-32481;
            end
    283   : begin
              real_value= 10783;
              imag_value=-30935;
            end
    284   : begin
              real_value= 16842;
              imag_value=-28100;
            end
    285   : begin
              real_value= 22199;
              imag_value=-24092;
            end
    286   : begin
              real_value= 26630;
              imag_value=-19081;
            end
    287   : begin
              real_value= 29950;
              imag_value=-13274;
            end
    288   : begin
              real_value= 32022;
              imag_value=-6915;
            end
    289   : begin
              real_value= 32759;
              imag_value=-267;
            end
    290   : begin
              real_value= 32131;
              imag_value=6390;
            end
    291   : begin
              real_value= 30163;
              imag_value=12784;
            end
    292   : begin
              real_value= 26938;
              imag_value=18644;
            end
    293   : begin
              real_value= 22589;
              imag_value=23726;
            end
    294   : begin
              real_value= 17299;
              imag_value=27820;
            end
    295   : begin
              real_value= 11289;
              imag_value=30755;
            end
    296   : begin
              real_value= 4806;
              imag_value=32407;
            end
    297   : begin
              real_value= -1874;
              imag_value=32707;
            end
    298   : begin
              real_value= -8477;
              imag_value=31645;
            end
    299   : begin
              real_value= -14728;
              imag_value=29263;
            end
    300   : begin
              real_value= -20365;
              imag_value=25661;
            end
    301   : begin
              real_value= -25154;
              imag_value=20988;
            end
    302   : begin
              real_value= -28892;
              imag_value=15442;
            end
    303   : begin
              real_value= -31426;
              imag_value=9253;
            end
    304   : begin
              real_value= -32651;
              imag_value=2676;
            end
    305   : begin
              real_value= -32515;
              imag_value=-4009;
            end
    306   : begin
              real_value= -31023;
              imag_value=-10529;
            end
    307   : begin
              real_value= -28236;
              imag_value=-16611;
            end
    308   : begin
              real_value= -24274;
              imag_value=-22001;
            end
    309   : begin
              real_value= -19299;
              imag_value=-26472;
            end
    310   : begin
              real_value= -13520;
              imag_value=-29841;
            end
    311   : begin
              real_value= -7177;
              imag_value=-31965;
            end
    312   : begin
              real_value= -535;
              imag_value=-32757;
            end
    313   : begin
              real_value= 6127;
              imag_value=-32183;
            end
    314   : begin
              real_value= 12537;
              imag_value=-30267;
            end
    315   : begin
              real_value= 18423;
              imag_value=-27090;
            end
    316   : begin
              real_value= 23541;
              imag_value=-22782;
            end
    317   : begin
              real_value= 27678;
              imag_value=-17525;
            end
    318   : begin
              real_value= 30661;
              imag_value=-11539;
            end
    319   : begin
              real_value= 32365;
              imag_value=-5071;
            end
    320   : begin
              real_value= 32721;
              imag_value=1606;
            end
    321   : begin
              real_value= 31713;
              imag_value=8219;
            end
    322   : begin
              real_value= 29382;
              imag_value=14489;
            end
    323   : begin
              real_value= 25826;
              imag_value=20154;
            end
    324   : begin
              real_value= 21194;
              imag_value=24981;
            end
    325   : begin
              real_value= 15678;
              imag_value=28766;
            end
    326   : begin
              real_value= 9508;
              imag_value=31351;
            end
    327   : begin
              real_value= 2942;
              imag_value=32629;
            end
    328   : begin
              real_value= -3742;
              imag_value=32547;
            end
    329   : begin
              real_value= -10275;
              imag_value=31107;
            end
    330   : begin
              real_value= -16380;
              imag_value=28371;
            end
    331   : begin
              real_value= -21801;
              imag_value=24453;
            end
    332   : begin
              real_value= -26314;
              imag_value=19515;
            end
    333   : begin
              real_value= -29729;
              imag_value=13764;
            end
    334   : begin
              real_value= -31905;
              imag_value=7438;
            end
    335   : begin
              real_value= -32750;
              imag_value=802;
            end
    336   : begin
              real_value= -32231;
              imag_value=-5864;
            end
    337   : begin
              real_value= -30369;
              imag_value=-12288;
            end
    338   : begin
              real_value= -27240;
              imag_value=-18200;
            end
    339   : begin
              real_value= -22974;
              imag_value=-23354;
            end
    340   : begin
              real_value= -17752;
              imag_value=-27534;
            end
    341   : begin
              real_value= -11790;
              imag_value=-30565;
            end
    342   : begin
              real_value= -5336;
              imag_value=-32323;
            end
    343   : begin
              real_value= 1338;
              imag_value=-32733;
            end
    344   : begin
              real_value= 7959;
              imag_value=-31779;
            end
    345   : begin
              real_value= 14248;
              imag_value=-29499;
            end
    346   : begin
              real_value= 19943;
              imag_value=-25990;
            end
    347   : begin
              real_value= 24806;
              imag_value=-21399;
            end
    348   : begin
              real_value= 28636;
              imag_value=-15914;
            end
    349   : begin
              real_value= 31271;
              imag_value=-9765;
            end
    350   : begin
              real_value= 32603;
              imag_value=-3210;
            end
    351   : begin
              real_value= 32575;
              imag_value=3476;
            end
    352   : begin
              real_value= 31191;
              imag_value=10021;
            end
    353   : begin
              real_value= 28506;
              imag_value=16148;
            end
    354   : begin
              real_value= 24630;
              imag_value=21600;
            end
    355   : begin
              real_value= 19729;
              imag_value=26152;
            end
    356   : begin
              real_value= 14006;
              imag_value=29615;
            end
    357   : begin
              real_value= 7699;
              imag_value=31843;
            end
    358   : begin
              real_value= 1070;
              imag_value=32743;
            end
    359   : begin
              real_value= -5599;
              imag_value=32278;
            end
    360   : begin
              real_value= -12039;
              imag_value=30468;
            end
    361   : begin
              real_value= -17977;
              imag_value=27387;
            end
    362   : begin
              real_value= -23165;
              imag_value=23165;
            end
    363   : begin
              real_value= -27387;
              imag_value=17977;
            end
    364   : begin
              real_value= -30468;
              imag_value=12039;
            end
    365   : begin
              real_value= -32278;
              imag_value=5599;
            end
    366   : begin
              real_value= -32743;
              imag_value=-1070;
            end
    367   : begin
              real_value= -31843;
              imag_value=-7699;
            end
    368   : begin
              real_value= -29615;
              imag_value=-14006;
            end
    369   : begin
              real_value= -26152;
              imag_value=-19729;
            end
    370   : begin
              real_value= -21600;
              imag_value=-24630;
            end
    371   : begin
              real_value= -16148;
              imag_value=-28506;
            end
    372   : begin
              real_value= -10021;
              imag_value=-31191;
            end
    373   : begin
              real_value= -3476;
              imag_value=-32575;
            end
    374   : begin
              real_value= 3210;
              imag_value=-32603;
            end
    375   : begin
              real_value= 9765;
              imag_value=-31271;
            end
    376   : begin
              real_value= 15914;
              imag_value=-28636;
            end
    377   : begin
              real_value= 21399;
              imag_value=-24806;
            end
    378   : begin
              real_value= 25990;
              imag_value=-19943;
            end
    379   : begin
              real_value= 29499;
              imag_value=-14248;
            end
    380   : begin
              real_value= 31779;
              imag_value=-7959;
            end
    381   : begin
              real_value= 32733;
              imag_value=-1338;
            end
    382   : begin
              real_value= 32323;
              imag_value=5336;
            end
    383   : begin
              real_value= 30565;
              imag_value=11790;
            end
    384   : begin
              real_value= 27534;
              imag_value=17752;
            end
    385   : begin
              real_value= 23354;
              imag_value=22974;
            end
    386   : begin
              real_value= 18200;
              imag_value=27240;
            end
    387   : begin
              real_value= 12288;
              imag_value=30369;
            end
    388   : begin
              real_value= 5864;
              imag_value=32231;
            end
    389   : begin
              real_value= -802;
              imag_value=32750;
            end
    390   : begin
              real_value= -7438;
              imag_value=31905;
            end
    391   : begin
              real_value= -13764;
              imag_value=29729;
            end
    392   : begin
              real_value= -19515;
              imag_value=26314;
            end
    393   : begin
              real_value= -24453;
              imag_value=21801;
            end
    394   : begin
              real_value= -28371;
              imag_value=16380;
            end
    395   : begin
              real_value= -31107;
              imag_value=10275;
            end
    396   : begin
              real_value= -32547;
              imag_value=3742;
            end
    397   : begin
              real_value= -32629;
              imag_value=-2942;
            end
    398   : begin
              real_value= -31351;
              imag_value=-9508;
            end
    399   : begin
              real_value= -28766;
              imag_value=-15678;
            end
    400   : begin
              real_value= -24981;
              imag_value=-21194;
            end
    401   : begin
              real_value= -20154;
              imag_value=-25826;
            end
    402   : begin
              real_value= -14489;
              imag_value=-29382;
            end
    403   : begin
              real_value= -8219;
              imag_value=-31713;
            end
    404   : begin
              real_value= -1606;
              imag_value=-32721;
            end
    405   : begin
              real_value= 5071;
              imag_value=-32365;
            end
    406   : begin
              real_value= 11539;
              imag_value=-30661;
            end
    407   : begin
              real_value= 17525;
              imag_value=-27678;
            end
    408   : begin
              real_value= 22782;
              imag_value=-23541;
            end
    409   : begin
              real_value= 27090;
              imag_value=-18423;
            end
    410   : begin
              real_value= 30267;
              imag_value=-12537;
            end
    411   : begin
              real_value= 32183;
              imag_value=-6127;
            end
    412   : begin
              real_value= 32757;
              imag_value=535;
            end
    413   : begin
              real_value= 31965;
              imag_value=7177;
            end
    414   : begin
              real_value= 29841;
              imag_value=13520;
            end
    415   : begin
              real_value= 26472;
              imag_value=19299;
            end
    416   : begin
              real_value= 22001;
              imag_value=24274;
            end
    417   : begin
              real_value= 16611;
              imag_value=28236;
            end
    418   : begin
              real_value= 10529;
              imag_value=31023;
            end
    419   : begin
              real_value= 4009;
              imag_value=32515;
            end
    420   : begin
              real_value= -2676;
              imag_value=32651;
            end
    421   : begin
              real_value= -9253;
              imag_value=31426;
            end
    422   : begin
              real_value= -15442;
              imag_value=28892;
            end
    423   : begin
              real_value= -20988;
              imag_value=25154;
            end
    424   : begin
              real_value= -25661;
              imag_value=20365;
            end
    425   : begin
              real_value= -29263;
              imag_value=14728;
            end
    426   : begin
              real_value= -31645;
              imag_value=8477;
            end
    427   : begin
              real_value= -32707;
              imag_value=1874;
            end
    428   : begin
              real_value= -32407;
              imag_value=-4806;
            end
    429   : begin
              real_value= -30755;
              imag_value=-11289;
            end
    430   : begin
              real_value= -27820;
              imag_value=-17299;
            end
    431   : begin
              real_value= -23726;
              imag_value=-22589;
            end
    432   : begin
              real_value= -18644;
              imag_value=-26938;
            end
    433   : begin
              real_value= -12784;
              imag_value=-30163;
            end
    434   : begin
              real_value= -6390;
              imag_value=-32131;
            end
    435   : begin
              real_value= 267;
              imag_value=-32759;
            end
    436   : begin
              real_value= 6915;
              imag_value=-32022;
            end
    437   : begin
              real_value= 13274;
              imag_value=-29950;
            end
    438   : begin
              real_value= 19081;
              imag_value=-26630;
            end
    439   : begin
              real_value= 24092;
              imag_value=-22199;
            end
    440   : begin
              real_value= 28100;
              imag_value=-16842;
            end
    441   : begin
              real_value= 30935;
              imag_value=-10783;
            end
    442   : begin
              real_value= 32481;
              imag_value=-4275;
            end
    443   : begin
              real_value= 32673;
              imag_value=2408;
            end
    444   : begin
              real_value= 31501;
              imag_value=8995;
            end
    445   : begin
              real_value= 29017;
              imag_value=15206;
            end
    446   : begin
              real_value= 25324;
              imag_value=20783;
            end
    447   : begin
              real_value= 20575;
              imag_value=25494;
            end
    448   : begin
              real_value= 14968;
              imag_value=29142;
            end
    449   : begin
              real_value= 8737;
              imag_value=31575;
            end
    450   : begin
              real_value= 2142;
              imag_value=32691;
            end
    451   : begin
              real_value= -4540;
              imag_value=32445;
            end
    452   : begin
              real_value= -11036;
              imag_value=30846;
            end
    453   : begin
              real_value= -17072;
              imag_value=27961;
            end
    454   : begin
              real_value= -22395;
              imag_value=23911;
            end
    455   : begin
              real_value= -26784;
              imag_value=18863;
            end
    456   : begin
              real_value= -30057;
              imag_value=13030;
            end
    457   : begin
              real_value= -32077;
              imag_value=6654;
            end
    458   : begin
              real_value= -32760;
              imag_value=0;
            end
    459   : begin
              real_value= -32077;
              imag_value=-6654;
            end
    460   : begin
              real_value= -30057;
              imag_value=-13030;
            end
    461   : begin
              real_value= -26784;
              imag_value=-18863;
            end
    462   : begin
              real_value= -22395;
              imag_value=-23911;
            end
    463   : begin
              real_value= -17072;
              imag_value=-27961;
            end
    464   : begin
              real_value= -11036;
              imag_value=-30846;
            end
    465   : begin
              real_value= -4540;
              imag_value=-32445;
            end
    466   : begin
              real_value= 2142;
              imag_value=-32691;
            end
    467   : begin
              real_value= 8737;
              imag_value=-31575;
            end
    468   : begin
              real_value= 14968;
              imag_value=-29142;
            end
    469   : begin
              real_value= 20575;
              imag_value=-25494;
            end
    470   : begin
              real_value= 25324;
              imag_value=-20783;
            end
    471   : begin
              real_value= 29017;
              imag_value=-15206;
            end
    472   : begin
              real_value= 31501;
              imag_value=-8995;
            end
    473   : begin
              real_value= 32673;
              imag_value=-2408;
            end
    474   : begin
              real_value= 32481;
              imag_value=4275;
            end
    475   : begin
              real_value= 30935;
              imag_value=10783;
            end
    476   : begin
              real_value= 28100;
              imag_value=16842;
            end
    477   : begin
              real_value= 24092;
              imag_value=22199;
            end
    478   : begin
              real_value= 19081;
              imag_value=26630;
            end
    479   : begin
              real_value= 13274;
              imag_value=29950;
            end
    480   : begin
              real_value= 6915;
              imag_value=32022;
            end
    481   : begin
              real_value= 267;
              imag_value=32759;
            end
    482   : begin
              real_value= -6390;
              imag_value=32131;
            end
    483   : begin
              real_value= -12784;
              imag_value=30163;
            end
    484   : begin
              real_value= -18644;
              imag_value=26938;
            end
    485   : begin
              real_value= -23726;
              imag_value=22589;
            end
    486   : begin
              real_value= -27820;
              imag_value=17299;
            end
    487   : begin
              real_value= -30755;
              imag_value=11289;
            end
    488   : begin
              real_value= -32407;
              imag_value=4806;
            end
    489   : begin
              real_value= -32707;
              imag_value=-1874;
            end
    490   : begin
              real_value= -31645;
              imag_value=-8477;
            end
    491   : begin
              real_value= -29263;
              imag_value=-14728;
            end
    492   : begin
              real_value= -25661;
              imag_value=-20365;
            end
    493   : begin
              real_value= -20988;
              imag_value=-25154;
            end
    494   : begin
              real_value= -15442;
              imag_value=-28892;
            end
    495   : begin
              real_value= -9253;
              imag_value=-31426;
            end
    496   : begin
              real_value= -2676;
              imag_value=-32651;
            end
    497   : begin
              real_value= 4009;
              imag_value=-32515;
            end
    498   : begin
              real_value= 10529;
              imag_value=-31023;
            end
    499   : begin
              real_value= 16611;
              imag_value=-28236;
            end
    500   : begin
              real_value= 22001;
              imag_value=-24274;
            end
    501   : begin
              real_value= 26472;
              imag_value=-19299;
            end
    502   : begin
              real_value= 29841;
              imag_value=-13520;
            end
    503   : begin
              real_value= 31965;
              imag_value=-7177;
            end
    504   : begin
              real_value= 32757;
              imag_value=-535;
            end
    505   : begin
              real_value= 32183;
              imag_value=6127;
            end
    506   : begin
              real_value= 30267;
              imag_value=12537;
            end
    507   : begin
              real_value= 27090;
              imag_value=18423;
            end
    508   : begin
              real_value= 22782;
              imag_value=23541;
            end
    509   : begin
              real_value= 17525;
              imag_value=27678;
            end
    510   : begin
              real_value= 11539;
              imag_value=30661;
            end
    511   : begin
              real_value= 5071;
              imag_value=32365;
            end
    512   : begin
              real_value= -1606;
              imag_value=32721;
            end
    513   : begin
              real_value= -8219;
              imag_value=31713;
            end
    514   : begin
              real_value= -14489;
              imag_value=29382;
            end
    515   : begin
              real_value= -20154;
              imag_value=25826;
            end
    516   : begin
              real_value= -24981;
              imag_value=21194;
            end
    517   : begin
              real_value= -28766;
              imag_value=15678;
            end
    518   : begin
              real_value= -31351;
              imag_value=9508;
            end
    519   : begin
              real_value= -32629;
              imag_value=2942;
            end
    520   : begin
              real_value= -32547;
              imag_value=-3742;
            end
    521   : begin
              real_value= -31107;
              imag_value=-10275;
            end
    522   : begin
              real_value= -28371;
              imag_value=-16380;
            end
    523   : begin
              real_value= -24453;
              imag_value=-21801;
            end
    524   : begin
              real_value= -19515;
              imag_value=-26314;
            end
    525   : begin
              real_value= -13764;
              imag_value=-29729;
            end
    526   : begin
              real_value= -7438;
              imag_value=-31905;
            end
    527   : begin
              real_value= -802;
              imag_value=-32750;
            end
    528   : begin
              real_value= 5864;
              imag_value=-32231;
            end
    529   : begin
              real_value= 12288;
              imag_value=-30369;
            end
    530   : begin
              real_value= 18200;
              imag_value=-27240;
            end
    531   : begin
              real_value= 23354;
              imag_value=-22974;
            end
    532   : begin
              real_value= 27534;
              imag_value=-17752;
            end
    533   : begin
              real_value= 30565;
              imag_value=-11790;
            end
    534   : begin
              real_value= 32323;
              imag_value=-5336;
            end
    535   : begin
              real_value= 32733;
              imag_value=1338;
            end
    536   : begin
              real_value= 31779;
              imag_value=7959;
            end
    537   : begin
              real_value= 29499;
              imag_value=14248;
            end
    538   : begin
              real_value= 25990;
              imag_value=19943;
            end
    539   : begin
              real_value= 21399;
              imag_value=24806;
            end
    540   : begin
              real_value= 15914;
              imag_value=28636;
            end
    541   : begin
              real_value= 9765;
              imag_value=31271;
            end
    542   : begin
              real_value= 3210;
              imag_value=32603;
            end
    543   : begin
              real_value= -3476;
              imag_value=32575;
            end
    544   : begin
              real_value= -10021;
              imag_value=31191;
            end
    545   : begin
              real_value= -16148;
              imag_value=28506;
            end
    546   : begin
              real_value= -21600;
              imag_value=24630;
            end
    547   : begin
              real_value= -26152;
              imag_value=19729;
            end
    548   : begin
              real_value= -29615;
              imag_value=14006;
            end
    549   : begin
              real_value= -31843;
              imag_value=7699;
            end
    550   : begin
              real_value= -32743;
              imag_value=1070;
            end
    551   : begin
              real_value= -32278;
              imag_value=-5599;
            end
    552   : begin
              real_value= -30468;
              imag_value=-12039;
            end
    553   : begin
              real_value= -27387;
              imag_value=-17977;
            end
    554   : begin
              real_value= -23165;
              imag_value=-23165;
            end
    555   : begin
              real_value= -17977;
              imag_value=-27387;
            end
    556   : begin
              real_value= -12039;
              imag_value=-30468;
            end
    557   : begin
              real_value= -5599;
              imag_value=-32278;
            end
    558   : begin
              real_value= 1070;
              imag_value=-32743;
            end
    559   : begin
              real_value= 7699;
              imag_value=-31843;
            end
    560   : begin
              real_value= 14006;
              imag_value=-29615;
            end
    561   : begin
              real_value= 19729;
              imag_value=-26152;
            end
    562   : begin
              real_value= 24630;
              imag_value=-21600;
            end
    563   : begin
              real_value= 28506;
              imag_value=-16148;
            end
    564   : begin
              real_value= 31191;
              imag_value=-10021;
            end
    565   : begin
              real_value= 32575;
              imag_value=-3476;
            end
    566   : begin
              real_value= 32603;
              imag_value=3210;
            end
    567   : begin
              real_value= 31271;
              imag_value=9765;
            end
    568   : begin
              real_value= 28636;
              imag_value=15914;
            end
    569   : begin
              real_value= 24806;
              imag_value=21399;
            end
    570   : begin
              real_value= 19943;
              imag_value=25990;
            end
    571   : begin
              real_value= 14248;
              imag_value=29499;
            end
    572   : begin
              real_value= 7959;
              imag_value=31779;
            end
    573   : begin
              real_value= 1338;
              imag_value=32733;
            end
    574   : begin
              real_value= -5336;
              imag_value=32323;
            end
    575   : begin
              real_value= -11790;
              imag_value=30565;
            end
    576   : begin
              real_value= -17752;
              imag_value=27534;
            end
    577   : begin
              real_value= -22974;
              imag_value=23354;
            end
    578   : begin
              real_value= -27240;
              imag_value=18200;
            end
    579   : begin
              real_value= -30369;
              imag_value=12288;
            end
    580   : begin
              real_value= -32231;
              imag_value=5864;
            end
    581   : begin
              real_value= -32750;
              imag_value=-802;
            end
    582   : begin
              real_value= -31905;
              imag_value=-7438;
            end
    583   : begin
              real_value= -29729;
              imag_value=-13764;
            end
    584   : begin
              real_value= -26314;
              imag_value=-19515;
            end
    585   : begin
              real_value= -21801;
              imag_value=-24453;
            end
    586   : begin
              real_value= -16380;
              imag_value=-28371;
            end
    587   : begin
              real_value= -10275;
              imag_value=-31107;
            end
    588   : begin
              real_value= -3742;
              imag_value=-32547;
            end
    589   : begin
              real_value= 2942;
              imag_value=-32629;
            end
    590   : begin
              real_value= 9508;
              imag_value=-31351;
            end
    591   : begin
              real_value= 15678;
              imag_value=-28766;
            end
    592   : begin
              real_value= 21194;
              imag_value=-24981;
            end
    593   : begin
              real_value= 25826;
              imag_value=-20154;
            end
    594   : begin
              real_value= 29382;
              imag_value=-14489;
            end
    595   : begin
              real_value= 31713;
              imag_value=-8219;
            end
    596   : begin
              real_value= 32721;
              imag_value=-1606;
            end
    597   : begin
              real_value= 32365;
              imag_value=5071;
            end
    598   : begin
              real_value= 30661;
              imag_value=11539;
            end
    599   : begin
              real_value= 27678;
              imag_value=17525;
            end
    600   : begin
              real_value= 23541;
              imag_value=22782;
            end
    601   : begin
              real_value= 18423;
              imag_value=27090;
            end
    602   : begin
              real_value= 12537;
              imag_value=30267;
            end
    603   : begin
              real_value= 6127;
              imag_value=32183;
            end
    604   : begin
              real_value= -535;
              imag_value=32757;
            end
    605   : begin
              real_value= -7177;
              imag_value=31965;
            end
    606   : begin
              real_value= -13520;
              imag_value=29841;
            end
    607   : begin
              real_value= -19299;
              imag_value=26472;
            end
    608   : begin
              real_value= -24274;
              imag_value=22001;
            end
    609   : begin
              real_value= -28236;
              imag_value=16611;
            end
    610   : begin
              real_value= -31023;
              imag_value=10529;
            end
    611   : begin
              real_value= -32515;
              imag_value=4009;
            end
    612   : begin
              real_value= -32651;
              imag_value=-2676;
            end
    613   : begin
              real_value= -31426;
              imag_value=-9253;
            end
    614   : begin
              real_value= -28892;
              imag_value=-15442;
            end
    615   : begin
              real_value= -25154;
              imag_value=-20988;
            end
    616   : begin
              real_value= -20365;
              imag_value=-25661;
            end
    617   : begin
              real_value= -14728;
              imag_value=-29263;
            end
    618   : begin
              real_value= -8477;
              imag_value=-31645;
            end
    619   : begin
              real_value= -1874;
              imag_value=-32707;
            end
    620   : begin
              real_value= 4806;
              imag_value=-32407;
            end
    621   : begin
              real_value= 11289;
              imag_value=-30755;
            end
    622   : begin
              real_value= 17299;
              imag_value=-27820;
            end
    623   : begin
              real_value= 22589;
              imag_value=-23726;
            end
    624   : begin
              real_value= 26938;
              imag_value=-18644;
            end
    625   : begin
              real_value= 30163;
              imag_value=-12784;
            end
    626   : begin
              real_value= 32131;
              imag_value=-6390;
            end
    627   : begin
              real_value= 32759;
              imag_value=267;
            end
    628   : begin
              real_value= 32022;
              imag_value=6915;
            end
    629   : begin
              real_value= 29950;
              imag_value=13274;
            end
    630   : begin
              real_value= 26630;
              imag_value=19081;
            end
    631   : begin
              real_value= 22199;
              imag_value=24092;
            end
    632   : begin
              real_value= 16842;
              imag_value=28100;
            end
    633   : begin
              real_value= 10783;
              imag_value=30935;
            end
    634   : begin
              real_value= 4275;
              imag_value=32481;
            end
    635   : begin
              real_value= -2408;
              imag_value=32673;
            end
    636   : begin
              real_value= -8995;
              imag_value=31501;
            end
    637   : begin
              real_value= -15206;
              imag_value=29017;
            end
    638   : begin
              real_value= -20783;
              imag_value=25324;
            end
    639   : begin
              real_value= -25494;
              imag_value=20575;
            end
    640   : begin
              real_value= -29142;
              imag_value=14968;
            end
    641   : begin
              real_value= -31575;
              imag_value=8737;
            end
    642   : begin
              real_value= -32691;
              imag_value=2142;
            end
    643   : begin
              real_value= -32445;
              imag_value=-4540;
            end
    644   : begin
              real_value= -30846;
              imag_value=-11036;
            end
    645   : begin
              real_value= -27961;
              imag_value=-17072;
            end
    646   : begin
              real_value= -23911;
              imag_value=-22395;
            end
    647   : begin
              real_value= -18863;
              imag_value=-26784;
            end
    648   : begin
              real_value= -13030;
              imag_value=-30057;
            end
    649   : begin
              real_value= -6654;
              imag_value=-32077;
            end
    650   : begin
              real_value= 0;
              imag_value=-32760;
            end
    651   : begin
              real_value= 6654;
              imag_value=-32077;
            end
    652   : begin
              real_value= 13030;
              imag_value=-30057;
            end
    653   : begin
              real_value= 18863;
              imag_value=-26784;
            end
    654   : begin
              real_value= 23911;
              imag_value=-22395;
            end
    655   : begin
              real_value= 27961;
              imag_value=-17072;
            end
    656   : begin
              real_value= 30846;
              imag_value=-11036;
            end
    657   : begin
              real_value= 32445;
              imag_value=-4540;
            end
    658   : begin
              real_value= 32691;
              imag_value=2142;
            end
    659   : begin
              real_value= 31575;
              imag_value=8737;
            end
    660   : begin
              real_value= 29142;
              imag_value=14968;
            end
    661   : begin
              real_value= 25494;
              imag_value=20575;
            end
    662   : begin
              real_value= 20783;
              imag_value=25324;
            end
    663   : begin
              real_value= 15206;
              imag_value=29017;
            end
    664   : begin
              real_value= 8995;
              imag_value=31501;
            end
    665   : begin
              real_value= 2408;
              imag_value=32673;
            end
    666   : begin
              real_value= -4275;
              imag_value=32481;
            end
    667   : begin
              real_value= -10783;
              imag_value=30935;
            end
    668   : begin
              real_value= -16842;
              imag_value=28100;
            end
    669   : begin
              real_value= -22199;
              imag_value=24092;
            end
    670   : begin
              real_value= -26630;
              imag_value=19081;
            end
    671   : begin
              real_value= -29950;
              imag_value=13274;
            end
    672   : begin
              real_value= -32022;
              imag_value=6915;
            end
    673   : begin
              real_value= -32759;
              imag_value=267;
            end
    674   : begin
              real_value= -32131;
              imag_value=-6390;
            end
    675   : begin
              real_value= -30163;
              imag_value=-12784;
            end
    676   : begin
              real_value= -26938;
              imag_value=-18644;
            end
    677   : begin
              real_value= -22589;
              imag_value=-23726;
            end
    678   : begin
              real_value= -17299;
              imag_value=-27820;
            end
    679   : begin
              real_value= -11289;
              imag_value=-30755;
            end
    680   : begin
              real_value= -4806;
              imag_value=-32407;
            end
    681   : begin
              real_value= 1874;
              imag_value=-32707;
            end
    682   : begin
              real_value= 8477;
              imag_value=-31645;
            end
    683   : begin
              real_value= 14728;
              imag_value=-29263;
            end
    684   : begin
              real_value= 20365;
              imag_value=-25661;
            end
    685   : begin
              real_value= 25154;
              imag_value=-20988;
            end
    686   : begin
              real_value= 28892;
              imag_value=-15442;
            end
    687   : begin
              real_value= 31426;
              imag_value=-9253;
            end
    688   : begin
              real_value= 32651;
              imag_value=-2676;
            end
    689   : begin
              real_value= 32515;
              imag_value=4009;
            end
    690   : begin
              real_value= 31023;
              imag_value=10529;
            end
    691   : begin
              real_value= 28236;
              imag_value=16611;
            end
    692   : begin
              real_value= 24274;
              imag_value=22001;
            end
    693   : begin
              real_value= 19299;
              imag_value=26472;
            end
    694   : begin
              real_value= 13520;
              imag_value=29841;
            end
    695   : begin
              real_value= 7177;
              imag_value=31965;
            end
    696   : begin
              real_value= 535;
              imag_value=32757;
            end
    697   : begin
              real_value= -6127;
              imag_value=32183;
            end
    698   : begin
              real_value= -12537;
              imag_value=30267;
            end
    699   : begin
              real_value= -18423;
              imag_value=27090;
            end
    700   : begin
              real_value= -23541;
              imag_value=22782;
            end
    701   : begin
              real_value= -27678;
              imag_value=17525;
            end
    702   : begin
              real_value= -30661;
              imag_value=11539;
            end
    703   : begin
              real_value= -32365;
              imag_value=5071;
            end
    704   : begin
              real_value= -32721;
              imag_value=-1606;
            end
    705   : begin
              real_value= -31713;
              imag_value=-8219;
            end
    706   : begin
              real_value= -29382;
              imag_value=-14489;
            end
    707   : begin
              real_value= -25826;
              imag_value=-20154;
            end
    708   : begin
              real_value= -21194;
              imag_value=-24981;
            end
    709   : begin
              real_value= -15678;
              imag_value=-28766;
            end
    710   : begin
              real_value= -9508;
              imag_value=-31351;
            end
    711   : begin
              real_value= -2942;
              imag_value=-32629;
            end
    712   : begin
              real_value= 3742;
              imag_value=-32547;
            end
    713   : begin
              real_value= 10275;
              imag_value=-31107;
            end
    714   : begin
              real_value= 16380;
              imag_value=-28371;
            end
    715   : begin
              real_value= 21801;
              imag_value=-24453;
            end
    716   : begin
              real_value= 26314;
              imag_value=-19515;
            end
    717   : begin
              real_value= 29729;
              imag_value=-13764;
            end
    718   : begin
              real_value= 31905;
              imag_value=-7438;
            end
    719   : begin
              real_value= 32750;
              imag_value=-802;
            end
    720   : begin
              real_value= 32231;
              imag_value=5864;
            end
    721   : begin
              real_value= 30369;
              imag_value=12288;
            end
    722   : begin
              real_value= 27240;
              imag_value=18200;
            end
    723   : begin
              real_value= 22974;
              imag_value=23354;
            end
    724   : begin
              real_value= 17752;
              imag_value=27534;
            end
    725   : begin
              real_value= 11790;
              imag_value=30565;
            end
    726   : begin
              real_value= 5336;
              imag_value=32323;
            end
    727   : begin
              real_value= -1338;
              imag_value=32733;
            end
    728   : begin
              real_value= -7959;
              imag_value=31779;
            end
    729   : begin
              real_value= -14248;
              imag_value=29499;
            end
    730   : begin
              real_value= -19943;
              imag_value=25990;
            end
    731   : begin
              real_value= -24806;
              imag_value=21399;
            end
    732   : begin
              real_value= -28636;
              imag_value=15914;
            end
    733   : begin
              real_value= -31271;
              imag_value=9765;
            end
    734   : begin
              real_value= -32603;
              imag_value=3210;
            end
    735   : begin
              real_value= -32575;
              imag_value=-3476;
            end
    736   : begin
              real_value= -31191;
              imag_value=-10021;
            end
    737   : begin
              real_value= -28506;
              imag_value=-16148;
            end
    738   : begin
              real_value= -24630;
              imag_value=-21600;
            end
    739   : begin
              real_value= -19729;
              imag_value=-26152;
            end
    740   : begin
              real_value= -14006;
              imag_value=-29615;
            end
    741   : begin
              real_value= -7699;
              imag_value=-31843;
            end
    742   : begin
              real_value= -1070;
              imag_value=-32743;
            end
    743   : begin
              real_value= 5599;
              imag_value=-32278;
            end
    744   : begin
              real_value= 12039;
              imag_value=-30468;
            end
    745   : begin
              real_value= 17977;
              imag_value=-27387;
            end
    746   : begin
              real_value= 23165;
              imag_value=-23165;
            end
    747   : begin
              real_value= 27387;
              imag_value=-17977;
            end
    748   : begin
              real_value= 30468;
              imag_value=-12039;
            end
    749   : begin
              real_value= 32278;
              imag_value=-5599;
            end
    750   : begin
              real_value= 32743;
              imag_value=1070;
            end
    751   : begin
              real_value= 31843;
              imag_value=7699;
            end
    752   : begin
              real_value= 29615;
              imag_value=14006;
            end
    753   : begin
              real_value= 26152;
              imag_value=19729;
            end
    754   : begin
              real_value= 21600;
              imag_value=24630;
            end
    755   : begin
              real_value= 16148;
              imag_value=28506;
            end
    756   : begin
              real_value= 10021;
              imag_value=31191;
            end
    757   : begin
              real_value= 3476;
              imag_value=32575;
            end
    758   : begin
              real_value= -3210;
              imag_value=32603;
            end
    759   : begin
              real_value= -9765;
              imag_value=31271;
            end
    760   : begin
              real_value= -15914;
              imag_value=28636;
            end
    761   : begin
              real_value= -21399;
              imag_value=24806;
            end
    762   : begin
              real_value= -25990;
              imag_value=19943;
            end
    763   : begin
              real_value= -29499;
              imag_value=14248;
            end
    764   : begin
              real_value= -31779;
              imag_value=7959;
            end
    765   : begin
              real_value= -32733;
              imag_value=1338;
            end
    766   : begin
              real_value= -32323;
              imag_value=-5336;
            end
    767   : begin
              real_value= -30565;
              imag_value=-11790;
            end
    768   : begin
              real_value= -27534;
              imag_value=-17752;
            end
    769   : begin
              real_value= -23354;
              imag_value=-22974;
            end
    770   : begin
              real_value= -18200;
              imag_value=-27240;
            end
    771   : begin
              real_value= -12288;
              imag_value=-30369;
            end
    772   : begin
              real_value= -5864;
              imag_value=-32231;
            end
    773   : begin
              real_value= 802;
              imag_value=-32750;
            end
    774   : begin
              real_value= 7438;
              imag_value=-31905;
            end
    775   : begin
              real_value= 13764;
              imag_value=-29729;
            end
    776   : begin
              real_value= 19515;
              imag_value=-26314;
            end
    777   : begin
              real_value= 24453;
              imag_value=-21801;
            end
    778   : begin
              real_value= 28371;
              imag_value=-16380;
            end
    779   : begin
              real_value= 31107;
              imag_value=-10275;
            end
    780   : begin
              real_value= 32547;
              imag_value=-3742;
            end
    781   : begin
              real_value= 32629;
              imag_value=2942;
            end
    782   : begin
              real_value= 31351;
              imag_value=9508;
            end
    783   : begin
              real_value= 28766;
              imag_value=15678;
            end
    784   : begin
              real_value= 24981;
              imag_value=21194;
            end
    785   : begin
              real_value= 20154;
              imag_value=25826;
            end
    786   : begin
              real_value= 14489;
              imag_value=29382;
            end
    787   : begin
              real_value= 8219;
              imag_value=31713;
            end
    788   : begin
              real_value= 1606;
              imag_value=32721;
            end
    789   : begin
              real_value= -5071;
              imag_value=32365;
            end
    790   : begin
              real_value= -11539;
              imag_value=30661;
            end
    791   : begin
              real_value= -17525;
              imag_value=27678;
            end
    792   : begin
              real_value= -22782;
              imag_value=23541;
            end
    793   : begin
              real_value= -27090;
              imag_value=18423;
            end
    794   : begin
              real_value= -30267;
              imag_value=12537;
            end
    795   : begin
              real_value= -32183;
              imag_value=6127;
            end
    796   : begin
              real_value= -32757;
              imag_value=-535;
            end
    797   : begin
              real_value= -31965;
              imag_value=-7177;
            end
    798   : begin
              real_value= -29841;
              imag_value=-13520;
            end
    799   : begin
              real_value= -26472;
              imag_value=-19299;
            end
    800   : begin
              real_value= -22001;
              imag_value=-24274;
            end
    801   : begin
              real_value= -16611;
              imag_value=-28236;
            end
    802   : begin
              real_value= -10529;
              imag_value=-31023;
            end
    803   : begin
              real_value= -4009;
              imag_value=-32515;
            end
    804   : begin
              real_value= 2676;
              imag_value=-32651;
            end
    805   : begin
              real_value= 9253;
              imag_value=-31426;
            end
    806   : begin
              real_value= 15442;
              imag_value=-28892;
            end
    807   : begin
              real_value= 20988;
              imag_value=-25154;
            end
    808   : begin
              real_value= 25661;
              imag_value=-20365;
            end
    809   : begin
              real_value= 29263;
              imag_value=-14728;
            end
    810   : begin
              real_value= 31645;
              imag_value=-8477;
            end
    811   : begin
              real_value= 32707;
              imag_value=-1874;
            end
    812   : begin
              real_value= 32407;
              imag_value=4806;
            end
    813   : begin
              real_value= 30755;
              imag_value=11289;
            end
    814   : begin
              real_value= 27820;
              imag_value=17299;
            end
    815   : begin
              real_value= 23726;
              imag_value=22589;
            end
    816   : begin
              real_value= 18644;
              imag_value=26938;
            end
    817   : begin
              real_value= 12784;
              imag_value=30163;
            end
    818   : begin
              real_value= 6390;
              imag_value=32131;
            end
    819   : begin
              real_value= -267;
              imag_value=32759;
            end
    820   : begin
              real_value= -6915;
              imag_value=32022;
            end
    821   : begin
              real_value= -13274;
              imag_value=29950;
            end
    822   : begin
              real_value= -19081;
              imag_value=26630;
            end
    823   : begin
              real_value= -24092;
              imag_value=22199;
            end
    824   : begin
              real_value= -28100;
              imag_value=16842;
            end
    825   : begin
              real_value= -30935;
              imag_value=10783;
            end
    826   : begin
              real_value= -32481;
              imag_value=4275;
            end
    827   : begin
              real_value= -32673;
              imag_value=-2408;
            end
    828   : begin
              real_value= -31501;
              imag_value=-8995;
            end
    829   : begin
              real_value= -29017;
              imag_value=-15206;
            end
    830   : begin
              real_value= -25324;
              imag_value=-20783;
            end
    831   : begin
              real_value= -20575;
              imag_value=-25494;
            end
    832   : begin
              real_value= -14968;
              imag_value=-29142;
            end
    833   : begin
              real_value= -8737;
              imag_value=-31575;
            end
    834   : begin
              real_value= -2142;
              imag_value=-32691;
            end
    835   : begin
              real_value= 4540;
              imag_value=-32445;
            end
    836   : begin
              real_value= 11036;
              imag_value=-30846;
            end
    837   : begin
              real_value= 17072;
              imag_value=-27961;
            end
    838   : begin
              real_value= 22395;
              imag_value=-23911;
            end
    839   : begin
              real_value= 26784;
              imag_value=-18863;
            end
    840   : begin
              real_value= 30057;
              imag_value=-13030;
            end
    841   : begin
              real_value= 32077;
              imag_value=-6654;
            end
    842   : begin
              real_value= 32760;
              imag_value=0;
            end
    843   : begin
              real_value= 32077;
              imag_value=6654;
            end
    844   : begin
              real_value= 30057;
              imag_value=13030;
            end
    845   : begin
              real_value= 26784;
              imag_value=18863;
            end
    846   : begin
              real_value= 22395;
              imag_value=23911;
            end
    847   : begin
              real_value= 17072;
              imag_value=27961;
            end
    848   : begin
              real_value= 11036;
              imag_value=30846;
            end
    849   : begin
              real_value= 4540;
              imag_value=32445;
            end
    850   : begin
              real_value= -2142;
              imag_value=32691;
            end
    851   : begin
              real_value= -8737;
              imag_value=31575;
            end
    852   : begin
              real_value= -14968;
              imag_value=29142;
            end
    853   : begin
              real_value= -20575;
              imag_value=25494;
            end
    854   : begin
              real_value= -25324;
              imag_value=20783;
            end
    855   : begin
              real_value= -29017;
              imag_value=15206;
            end
    856   : begin
              real_value= -31501;
              imag_value=8995;
            end
    857   : begin
              real_value= -32673;
              imag_value=2408;
            end
    858   : begin
              real_value= -32481;
              imag_value=-4275;
            end
    859   : begin
              real_value= -30935;
              imag_value=-10783;
            end
    860   : begin
              real_value= -28100;
              imag_value=-16842;
            end
    861   : begin
              real_value= -24092;
              imag_value=-22199;
            end
    862   : begin
              real_value= -19081;
              imag_value=-26630;
            end
    863   : begin
              real_value= -13274;
              imag_value=-29950;
            end
    864   : begin
              real_value= -6915;
              imag_value=-32022;
            end
    865   : begin
              real_value= -267;
              imag_value=-32759;
            end
    866   : begin
              real_value= 6390;
              imag_value=-32131;
            end
    867   : begin
              real_value= 12784;
              imag_value=-30163;
            end
    868   : begin
              real_value= 18644;
              imag_value=-26938;
            end
    869   : begin
              real_value= 23726;
              imag_value=-22589;
            end
    870   : begin
              real_value= 27820;
              imag_value=-17299;
            end
    871   : begin
              real_value= 30755;
              imag_value=-11289;
            end
    872   : begin
              real_value= 32407;
              imag_value=-4806;
            end
    873   : begin
              real_value= 32707;
              imag_value=1874;
            end
    874   : begin
              real_value= 31645;
              imag_value=8477;
            end
    875   : begin
              real_value= 29263;
              imag_value=14728;
            end
    876   : begin
              real_value= 25661;
              imag_value=20365;
            end
    877   : begin
              real_value= 20988;
              imag_value=25154;
            end
    878   : begin
              real_value= 15442;
              imag_value=28892;
            end
    879   : begin
              real_value= 9253;
              imag_value=31426;
            end
    880   : begin
              real_value= 2676;
              imag_value=32651;
            end
    881   : begin
              real_value= -4009;
              imag_value=32515;
            end
    882   : begin
              real_value= -10529;
              imag_value=31023;
            end
    883   : begin
              real_value= -16611;
              imag_value=28236;
            end
    884   : begin
              real_value= -22001;
              imag_value=24274;
            end
    885   : begin
              real_value= -26472;
              imag_value=19299;
            end
    886   : begin
              real_value= -29841;
              imag_value=13520;
            end
    887   : begin
              real_value= -31965;
              imag_value=7177;
            end
    888   : begin
              real_value= -32757;
              imag_value=535;
            end
    889   : begin
              real_value= -32183;
              imag_value=-6127;
            end
    890   : begin
              real_value= -30267;
              imag_value=-12537;
            end
    891   : begin
              real_value= -27090;
              imag_value=-18423;
            end
    892   : begin
              real_value= -22782;
              imag_value=-23541;
            end
    893   : begin
              real_value= -17525;
              imag_value=-27678;
            end
    894   : begin
              real_value= -11539;
              imag_value=-30661;
            end
    895   : begin
              real_value= -5071;
              imag_value=-32365;
            end
    896   : begin
              real_value= 1606;
              imag_value=-32721;
            end
    897   : begin
              real_value= 8219;
              imag_value=-31713;
            end
    898   : begin
              real_value= 14489;
              imag_value=-29382;
            end
    899   : begin
              real_value= 20154;
              imag_value=-25826;
            end
    900   : begin
              real_value= 24981;
              imag_value=-21194;
            end
    901   : begin
              real_value= 28766;
              imag_value=-15678;
            end
    902   : begin
              real_value= 31351;
              imag_value=-9508;
            end
    903   : begin
              real_value= 32629;
              imag_value=-2942;
            end
    904   : begin
              real_value= 32547;
              imag_value=3742;
            end
    905   : begin
              real_value= 31107;
              imag_value=10275;
            end
    906   : begin
              real_value= 28371;
              imag_value=16380;
            end
    907   : begin
              real_value= 24453;
              imag_value=21801;
            end
    908   : begin
              real_value= 19515;
              imag_value=26314;
            end
    909   : begin
              real_value= 13764;
              imag_value=29729;
            end
    910   : begin
              real_value= 7438;
              imag_value=31905;
            end
    911   : begin
              real_value= 802;
              imag_value=32750;
            end
    912   : begin
              real_value= -5864;
              imag_value=32231;
            end
    913   : begin
              real_value= -12288;
              imag_value=30369;
            end
    914   : begin
              real_value= -18200;
              imag_value=27240;
            end
    915   : begin
              real_value= -23354;
              imag_value=22974;
            end
    916   : begin
              real_value= -27534;
              imag_value=17752;
            end
    917   : begin
              real_value= -30565;
              imag_value=11790;
            end
    918   : begin
              real_value= -32323;
              imag_value=5336;
            end
    919   : begin
              real_value= -32733;
              imag_value=-1338;
            end
    920   : begin
              real_value= -31779;
              imag_value=-7959;
            end
    921   : begin
              real_value= -29499;
              imag_value=-14248;
            end
    922   : begin
              real_value= -25990;
              imag_value=-19943;
            end
    923   : begin
              real_value= -21399;
              imag_value=-24806;
            end
    924   : begin
              real_value= -15914;
              imag_value=-28636;
            end
    925   : begin
              real_value= -9765;
              imag_value=-31271;
            end
    926   : begin
              real_value= -3210;
              imag_value=-32603;
            end
    927   : begin
              real_value= 3476;
              imag_value=-32575;
            end
    928   : begin
              real_value= 10021;
              imag_value=-31191;
            end
    929   : begin
              real_value= 16148;
              imag_value=-28506;
            end
    930   : begin
              real_value= 21600;
              imag_value=-24630;
            end
    931   : begin
              real_value= 26152;
              imag_value=-19729;
            end
    932   : begin
              real_value= 29615;
              imag_value=-14006;
            end
    933   : begin
              real_value= 31843;
              imag_value=-7699;
            end
    934   : begin
              real_value= 32743;
              imag_value=-1070;
            end
    935   : begin
              real_value= 32278;
              imag_value=5599;
            end
    936   : begin
              real_value= 30468;
              imag_value=12039;
            end
    937   : begin
              real_value= 27387;
              imag_value=17977;
            end
    938   : begin
              real_value= 23165;
              imag_value=23165;
            end
    939   : begin
              real_value= 17977;
              imag_value=27387;
            end
    940   : begin
              real_value= 12039;
              imag_value=30468;
            end
    941   : begin
              real_value= 5599;
              imag_value=32278;
            end
    942   : begin
              real_value= -1070;
              imag_value=32743;
            end
    943   : begin
              real_value= -7699;
              imag_value=31843;
            end
    944   : begin
              real_value= -14006;
              imag_value=29615;
            end
    945   : begin
              real_value= -19729;
              imag_value=26152;
            end
    946   : begin
              real_value= -24630;
              imag_value=21600;
            end
    947   : begin
              real_value= -28506;
              imag_value=16148;
            end
    948   : begin
              real_value= -31191;
              imag_value=10021;
            end
    949   : begin
              real_value= -32575;
              imag_value=3476;
            end
    950   : begin
              real_value= -32603;
              imag_value=-3210;
            end
    951   : begin
              real_value= -31271;
              imag_value=-9765;
            end
    952   : begin
              real_value= -28636;
              imag_value=-15914;
            end
    953   : begin
              real_value= -24806;
              imag_value=-21399;
            end
    954   : begin
              real_value= -19943;
              imag_value=-25990;
            end
    955   : begin
              real_value= -14248;
              imag_value=-29499;
            end
    956   : begin
              real_value= -7959;
              imag_value=-31779;
            end
    957   : begin
              real_value= -1338;
              imag_value=-32733;
            end
    958   : begin
              real_value= 5336;
              imag_value=-32323;
            end
    959   : begin
              real_value= 11790;
              imag_value=-30565;
            end
    960   : begin
              real_value= 17752;
              imag_value=-27534;
            end
    961   : begin
              real_value= 22974;
              imag_value=-23354;
            end
    962   : begin
              real_value= 27240;
              imag_value=-18200;
            end
    963   : begin
              real_value= 30369;
              imag_value=-12288;
            end
    964   : begin
              real_value= 32231;
              imag_value=-5864;
            end
    965   : begin
              real_value= 32750;
              imag_value=802;
            end
    966   : begin
              real_value= 31905;
              imag_value=7438;
            end
    967   : begin
              real_value= 29729;
              imag_value=13764;
            end
    968   : begin
              real_value= 26314;
              imag_value=19515;
            end
    969   : begin
              real_value= 21801;
              imag_value=24453;
            end
    970   : begin
              real_value= 16380;
              imag_value=28371;
            end
    971   : begin
              real_value= 10275;
              imag_value=31107;
            end
    972   : begin
              real_value= 3742;
              imag_value=32547;
            end
    973   : begin
              real_value= -2942;
              imag_value=32629;
            end
    974   : begin
              real_value= -9508;
              imag_value=31351;
            end
    975   : begin
              real_value= -15678;
              imag_value=28766;
            end
    976   : begin
              real_value= -21194;
              imag_value=24981;
            end
    977   : begin
              real_value= -25826;
              imag_value=20154;
            end
    978   : begin
              real_value= -29382;
              imag_value=14489;
            end
    979   : begin
              real_value= -31713;
              imag_value=8219;
            end
    980   : begin
              real_value= -32721;
              imag_value=1606;
            end
    981   : begin
              real_value= -32365;
              imag_value=-5071;
            end
    982   : begin
              real_value= -30661;
              imag_value=-11539;
            end
    983   : begin
              real_value= -27678;
              imag_value=-17525;
            end
    984   : begin
              real_value= -23541;
              imag_value=-22782;
            end
    985   : begin
              real_value= -18423;
              imag_value=-27090;
            end
    986   : begin
              real_value= -12537;
              imag_value=-30267;
            end
    987   : begin
              real_value= -6127;
              imag_value=-32183;
            end
    988   : begin
              real_value= 535;
              imag_value=-32757;
            end
    989   : begin
              real_value= 7177;
              imag_value=-31965;
            end
    990   : begin
              real_value= 13520;
              imag_value=-29841;
            end
    991   : begin
              real_value= 19299;
              imag_value=-26472;
            end
    992   : begin
              real_value= 24274;
              imag_value=-22001;
            end
    993   : begin
              real_value= 28236;
              imag_value=-16611;
            end
    994   : begin
              real_value= 31023;
              imag_value=-10529;
            end
    995   : begin
              real_value= 32515;
              imag_value=-4009;
            end
    996   : begin
              real_value= 32651;
              imag_value=2676;
            end
    997   : begin
              real_value= 31426;
              imag_value=9253;
            end
    998   : begin
              real_value= 28892;
              imag_value=15442;
            end
    999   : begin
              real_value= 25154;
              imag_value=20988;
            end
    1000   : begin
              real_value= 20365;
              imag_value=25661;
            end
    1001  : begin
              real_value= 14728;
              imag_value=29263;
            end
    1002  : begin
              real_value= 8477;
              imag_value=31645;
            end
    1003  : begin
              real_value= 1874;
              imag_value=32707;
            end
    1004  : begin
              real_value= -4806;
              imag_value=32407;
            end
    1005  : begin
              real_value= -11289;
              imag_value=30755;
            end
    1006  : begin
              real_value= -17299;
              imag_value=27820;
            end
    1007  : begin
              real_value= -22589;
              imag_value=23726;
            end
    1008  : begin
              real_value= -26938;
              imag_value=18644;
            end
    1009  : begin
              real_value= -30163;
              imag_value=12784;
            end
    1010  : begin
              real_value= -32131;
              imag_value=6390;
            end
    1011  : begin
              real_value= -32759;
              imag_value=-267;
            end
    1012  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    1013  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    1014  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    1015  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    1016  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    1017  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    1018  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    1019  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    1020  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    1021  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    1022  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    1023  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    1024  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    1025  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    1026  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    1027  : begin
              real_value= 32445;
              imag_value=4540;
            end
    1028  : begin
              real_value= 30846;
              imag_value=11036;
            end
    1029  : begin
              real_value= 27961;
              imag_value=17072;
            end
    1030  : begin
              real_value= 23911;
              imag_value=22395;
            end
    1031  : begin
              real_value= 18863;
              imag_value=26784;
            end
    1032  : begin
              real_value= 13030;
              imag_value=30057;
            end
    1033  : begin
              real_value= 6654;
              imag_value=32077;
            end
    1034  : begin
              real_value= 0;
              imag_value=32760;
            end
    1035  : begin
              real_value= -6654;
              imag_value=32077;
            end
    1036  : begin
              real_value= -13030;
              imag_value=30057;
            end
    1037  : begin
              real_value= -18863;
              imag_value=26784;
            end
    1038  : begin
              real_value= -23911;
              imag_value=22395;
            end
    1039  : begin
              real_value= -27961;
              imag_value=17072;
            end
    1040  : begin
              real_value= -30846;
              imag_value=11036;
            end
    1041  : begin
              real_value= -32445;
              imag_value=4540;
            end
    1042  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    1043  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    1044  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    1045  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    1046  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    1047  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    1048  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    1049  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    1050  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    1051  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    1052  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    1053  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    1054  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    1055  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    1056  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    1057  : begin
              real_value= 32759;
              imag_value=-267;
            end
    1058  : begin
              real_value= 32131;
              imag_value=6390;
            end
    1059  : begin
              real_value= 30163;
              imag_value=12784;
            end
    1060  : begin
              real_value= 26938;
              imag_value=18644;
            end
    1061  : begin
              real_value= 22589;
              imag_value=23726;
            end
    1062  : begin
              real_value= 17299;
              imag_value=27820;
            end
    1063  : begin
              real_value= 11289;
              imag_value=30755;
            end
    1064  : begin
              real_value= 4806;
              imag_value=32407;
            end
    1065  : begin
              real_value= -1874;
              imag_value=32707;
            end
    1066  : begin
              real_value= -8477;
              imag_value=31645;
            end
    1067  : begin
              real_value= -14728;
              imag_value=29263;
            end
    1068  : begin
              real_value= -20365;
              imag_value=25661;
            end
    1069  : begin
              real_value= -25154;
              imag_value=20988;
            end
    1070  : begin
              real_value= -28892;
              imag_value=15442;
            end
    1071  : begin
              real_value= -31426;
              imag_value=9253;
            end
    1072  : begin
              real_value= -32651;
              imag_value=2676;
            end
    1073  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    1074  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    1075  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    1076  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    1077  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    1078  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    1079  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    1080  : begin
              real_value= -535;
              imag_value=-32757;
            end
    1081  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    1082  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    1083  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    1084  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    1085  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    1086  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    1087  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    1088  : begin
              real_value= 32721;
              imag_value=1606;
            end
    1089  : begin
              real_value= 31713;
              imag_value=8219;
            end
    1090  : begin
              real_value= 29382;
              imag_value=14489;
            end
    1091  : begin
              real_value= 25826;
              imag_value=20154;
            end
    1092  : begin
              real_value= 21194;
              imag_value=24981;
            end
    1093  : begin
              real_value= 15678;
              imag_value=28766;
            end
    1094  : begin
              real_value= 9508;
              imag_value=31351;
            end
    1095  : begin
              real_value= 2942;
              imag_value=32629;
            end
    1096  : begin
              real_value= -3742;
              imag_value=32547;
            end
    1097  : begin
              real_value= -10275;
              imag_value=31107;
            end
    1098  : begin
              real_value= -16380;
              imag_value=28371;
            end
    1099  : begin
              real_value= -21801;
              imag_value=24453;
            end
    1100  : begin
              real_value= -26314;
              imag_value=19515;
            end
    1101  : begin
              real_value= -29729;
              imag_value=13764;
            end
    1102  : begin
              real_value= -31905;
              imag_value=7438;
            end
    1103  : begin
              real_value= -32750;
              imag_value=802;
            end
    1104  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    1105  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    1106  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    1107  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    1108  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    1109  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    1110  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    1111  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    1112  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    1113  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    1114  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    1115  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    1116  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    1117  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    1118  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    1119  : begin
              real_value= 32575;
              imag_value=3476;
            end
    1120  : begin
              real_value= 31191;
              imag_value=10021;
            end
    1121  : begin
              real_value= 28506;
              imag_value=16148;
            end
    1122  : begin
              real_value= 24630;
              imag_value=21600;
            end
    1123  : begin
              real_value= 19729;
              imag_value=26152;
            end
    1124  : begin
              real_value= 14006;
              imag_value=29615;
            end
    1125  : begin
              real_value= 7699;
              imag_value=31843;
            end
    1126  : begin
              real_value= 1070;
              imag_value=32743;
            end
    1127  : begin
              real_value= -5599;
              imag_value=32278;
            end
    1128  : begin
              real_value= -12039;
              imag_value=30468;
            end
    1129  : begin
              real_value= -17977;
              imag_value=27387;
            end
    1130  : begin
              real_value= -23165;
              imag_value=23165;
            end
    1131  : begin
              real_value= -27387;
              imag_value=17977;
            end
    1132  : begin
              real_value= -30468;
              imag_value=12039;
            end
    1133  : begin
              real_value= -32278;
              imag_value=5599;
            end
    1134  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    1135  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    1136  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    1137  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    1138  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    1139  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    1140  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    1141  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    1142  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    1143  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    1144  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    1145  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    1146  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    1147  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    1148  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    1149  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    1150  : begin
              real_value= 32323;
              imag_value=5336;
            end
    1151  : begin
              real_value= 30565;
              imag_value=11790;
            end
    1152  : begin
              real_value= 27534;
              imag_value=17752;
            end
    1153  : begin
              real_value= 23354;
              imag_value=22974;
            end
    1154  : begin
              real_value= 18200;
              imag_value=27240;
            end
    1155  : begin
              real_value= 12288;
              imag_value=30369;
            end
    1156  : begin
              real_value= 5864;
              imag_value=32231;
            end
    1157  : begin
              real_value= -802;
              imag_value=32750;
            end
    1158  : begin
              real_value= -7438;
              imag_value=31905;
            end
    1159  : begin
              real_value= -13764;
              imag_value=29729;
            end
    1160  : begin
              real_value= -19515;
              imag_value=26314;
            end
    1161  : begin
              real_value= -24453;
              imag_value=21801;
            end
    1162  : begin
              real_value= -28371;
              imag_value=16380;
            end
    1163  : begin
              real_value= -31107;
              imag_value=10275;
            end
    1164  : begin
              real_value= -32547;
              imag_value=3742;
            end
    1165  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    1166  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    1167  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    1168  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    1169  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    1170  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    1171  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    1172  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    1173  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    1174  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    1175  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    1176  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    1177  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    1178  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    1179  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    1180  : begin
              real_value= 32757;
              imag_value=535;
            end
    1181  : begin
              real_value= 31965;
              imag_value=7177;
            end
    1182  : begin
              real_value= 29841;
              imag_value=13520;
            end
    1183  : begin
              real_value= 26472;
              imag_value=19299;
            end
    1184  : begin
              real_value= 22001;
              imag_value=24274;
            end
    1185  : begin
              real_value= 16611;
              imag_value=28236;
            end
    1186  : begin
              real_value= 10529;
              imag_value=31023;
            end
    1187  : begin
              real_value= 4009;
              imag_value=32515;
            end
    1188  : begin
              real_value= -2676;
              imag_value=32651;
            end
    1189  : begin
              real_value= -9253;
              imag_value=31426;
            end
    1190  : begin
              real_value= -15442;
              imag_value=28892;
            end
    1191  : begin
              real_value= -20988;
              imag_value=25154;
            end
    1192  : begin
              real_value= -25661;
              imag_value=20365;
            end
    1193  : begin
              real_value= -29263;
              imag_value=14728;
            end
    1194  : begin
              real_value= -31645;
              imag_value=8477;
            end
    1195  : begin
              real_value= -32707;
              imag_value=1874;
            end
    1196  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    1197  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    1198  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    1199  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    1200  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    1201  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    1202  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    1203  : begin
              real_value= 267;
              imag_value=-32759;
            end
    1204  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    1205  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    1206  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    1207  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    1208  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    1209  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    1210  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    1211  : begin
              real_value= 32673;
              imag_value=2408;
            end
    1212  : begin
              real_value= 31501;
              imag_value=8995;
            end
    1213  : begin
              real_value= 29017;
              imag_value=15206;
            end
    1214  : begin
              real_value= 25324;
              imag_value=20783;
            end
    1215  : begin
              real_value= 20575;
              imag_value=25494;
            end
    1216  : begin
              real_value= 14968;
              imag_value=29142;
            end
    1217  : begin
              real_value= 8737;
              imag_value=31575;
            end
    1218  : begin
              real_value= 2142;
              imag_value=32691;
            end
    1219  : begin
              real_value= -4540;
              imag_value=32445;
            end
    1220  : begin
              real_value= -11036;
              imag_value=30846;
            end
    1221  : begin
              real_value= -17072;
              imag_value=27961;
            end
    1222  : begin
              real_value= -22395;
              imag_value=23911;
            end
    1223  : begin
              real_value= -26784;
              imag_value=18863;
            end
    1224  : begin
              real_value= -30057;
              imag_value=13030;
            end
    1225  : begin
              real_value= -32077;
              imag_value=6654;
            end
    1226  : begin
              real_value= -32760;
              imag_value=0;
            end
    1227  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    1228  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    1229  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    1230  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    1231  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    1232  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    1233  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    1234  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    1235  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    1236  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    1237  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    1238  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    1239  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    1240  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    1241  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    1242  : begin
              real_value= 32481;
              imag_value=4275;
            end
    1243  : begin
              real_value= 30935;
              imag_value=10783;
            end
    1244  : begin
              real_value= 28100;
              imag_value=16842;
            end
    1245  : begin
              real_value= 24092;
              imag_value=22199;
            end
    1246  : begin
              real_value= 19081;
              imag_value=26630;
            end
    1247  : begin
              real_value= 13274;
              imag_value=29950;
            end
    1248  : begin
              real_value= 6915;
              imag_value=32022;
            end
    1249  : begin
              real_value= 267;
              imag_value=32759;
            end
    1250  : begin
              real_value= -6390;
              imag_value=32131;
            end
    1251  : begin
              real_value= -12784;
              imag_value=30163;
            end
    1252  : begin
              real_value= -18644;
              imag_value=26938;
            end
    1253  : begin
              real_value= -23726;
              imag_value=22589;
            end
    1254  : begin
              real_value= -27820;
              imag_value=17299;
            end
    1255  : begin
              real_value= -30755;
              imag_value=11289;
            end
    1256  : begin
              real_value= -32407;
              imag_value=4806;
            end
    1257  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    1258  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    1259  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    1260  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    1261  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    1262  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    1263  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    1264  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    1265  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    1266  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    1267  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    1268  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    1269  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    1270  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    1271  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    1272  : begin
              real_value= 32757;
              imag_value=-535;
            end
    1273  : begin
              real_value= 32183;
              imag_value=6127;
            end
    1274  : begin
              real_value= 30267;
              imag_value=12537;
            end
    1275  : begin
              real_value= 27090;
              imag_value=18423;
            end
    1276  : begin
              real_value= 22782;
              imag_value=23541;
            end
    1277  : begin
              real_value= 17525;
              imag_value=27678;
            end
    1278  : begin
              real_value= 11539;
              imag_value=30661;
            end
    1279  : begin
              real_value= 5071;
              imag_value=32365;
            end
    1280  : begin
              real_value= -1606;
              imag_value=32721;
            end
    1281  : begin
              real_value= -8219;
              imag_value=31713;
            end
    1282  : begin
              real_value= -14489;
              imag_value=29382;
            end
    1283  : begin
              real_value= -20154;
              imag_value=25826;
            end
    1284  : begin
              real_value= -24981;
              imag_value=21194;
            end
    1285  : begin
              real_value= -28766;
              imag_value=15678;
            end
    1286  : begin
              real_value= -31351;
              imag_value=9508;
            end
    1287  : begin
              real_value= -32629;
              imag_value=2942;
            end
    1288  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    1289  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    1290  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    1291  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    1292  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    1293  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    1294  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    1295  : begin
              real_value= -802;
              imag_value=-32750;
            end
    1296  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    1297  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    1298  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    1299  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    1300  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    1301  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    1302  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    1303  : begin
              real_value= 32733;
              imag_value=1338;
            end
    1304  : begin
              real_value= 31779;
              imag_value=7959;
            end
    1305  : begin
              real_value= 29499;
              imag_value=14248;
            end
    1306  : begin
              real_value= 25990;
              imag_value=19943;
            end
    1307  : begin
              real_value= 21399;
              imag_value=24806;
            end
    1308  : begin
              real_value= 15914;
              imag_value=28636;
            end
    1309  : begin
              real_value= 9765;
              imag_value=31271;
            end
    1310  : begin
              real_value= 3210;
              imag_value=32603;
            end
    1311  : begin
              real_value= -3476;
              imag_value=32575;
            end
    1312  : begin
              real_value= -10021;
              imag_value=31191;
            end
    1313  : begin
              real_value= -16148;
              imag_value=28506;
            end
    1314  : begin
              real_value= -21600;
              imag_value=24630;
            end
    1315  : begin
              real_value= -26152;
              imag_value=19729;
            end
    1316  : begin
              real_value= -29615;
              imag_value=14006;
            end
    1317  : begin
              real_value= -31843;
              imag_value=7699;
            end
    1318  : begin
              real_value= -32743;
              imag_value=1070;
            end
    1319  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    1320  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    1321  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    1322  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    1323  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    1324  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    1325  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    1326  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    1327  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    1328  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    1329  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    1330  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    1331  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    1332  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    1333  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    1334  : begin
              real_value= 32603;
              imag_value=3210;
            end
    1335  : begin
              real_value= 31271;
              imag_value=9765;
            end
    1336  : begin
              real_value= 28636;
              imag_value=15914;
            end
    1337  : begin
              real_value= 24806;
              imag_value=21399;
            end
    1338  : begin
              real_value= 19943;
              imag_value=25990;
            end
    1339  : begin
              real_value= 14248;
              imag_value=29499;
            end
    1340  : begin
              real_value= 7959;
              imag_value=31779;
            end
    1341  : begin
              real_value= 1338;
              imag_value=32733;
            end
    1342  : begin
              real_value= -5336;
              imag_value=32323;
            end
    1343  : begin
              real_value= -11790;
              imag_value=30565;
            end
    1344  : begin
              real_value= -17752;
              imag_value=27534;
            end
    1345  : begin
              real_value= -22974;
              imag_value=23354;
            end
    1346  : begin
              real_value= -27240;
              imag_value=18200;
            end
    1347  : begin
              real_value= -30369;
              imag_value=12288;
            end
    1348  : begin
              real_value= -32231;
              imag_value=5864;
            end
    1349  : begin
              real_value= -32750;
              imag_value=-802;
            end
    1350  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    1351  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    1352  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    1353  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    1354  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    1355  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    1356  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    1357  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    1358  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    1359  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    1360  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    1361  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    1362  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    1363  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    1364  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    1365  : begin
              real_value= 32365;
              imag_value=5071;
            end
    1366  : begin
              real_value= 30661;
              imag_value=11539;
            end
    1367  : begin
              real_value= 27678;
              imag_value=17525;
            end
    1368  : begin
              real_value= 23541;
              imag_value=22782;
            end
    1369  : begin
              real_value= 18423;
              imag_value=27090;
            end
    1370  : begin
              real_value= 12537;
              imag_value=30267;
            end
    1371  : begin
              real_value= 6127;
              imag_value=32183;
            end
    1372  : begin
              real_value= -535;
              imag_value=32757;
            end
    1373  : begin
              real_value= -7177;
              imag_value=31965;
            end
    1374  : begin
              real_value= -13520;
              imag_value=29841;
            end
    1375  : begin
              real_value= -19299;
              imag_value=26472;
            end
    1376  : begin
              real_value= -24274;
              imag_value=22001;
            end
    1377  : begin
              real_value= -28236;
              imag_value=16611;
            end
    1378  : begin
              real_value= -31023;
              imag_value=10529;
            end
    1379  : begin
              real_value= -32515;
              imag_value=4009;
            end
    1380  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    1381  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    1382  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    1383  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    1384  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    1385  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    1386  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    1387  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    1388  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    1389  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    1390  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    1391  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    1392  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    1393  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    1394  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    1395  : begin
              real_value= 32759;
              imag_value=267;
            end
    1396  : begin
              real_value= 32022;
              imag_value=6915;
            end
    1397  : begin
              real_value= 29950;
              imag_value=13274;
            end
    1398  : begin
              real_value= 26630;
              imag_value=19081;
            end
    1399  : begin
              real_value= 22199;
              imag_value=24092;
            end
    1400  : begin
              real_value= 16842;
              imag_value=28100;
            end
    1401  : begin
              real_value= 10783;
              imag_value=30935;
            end
    1402  : begin
              real_value= 4275;
              imag_value=32481;
            end
    1403  : begin
              real_value= -2408;
              imag_value=32673;
            end
    1404  : begin
              real_value= -8995;
              imag_value=31501;
            end
    1405  : begin
              real_value= -15206;
              imag_value=29017;
            end
    1406  : begin
              real_value= -20783;
              imag_value=25324;
            end
    1407  : begin
              real_value= -25494;
              imag_value=20575;
            end
    1408  : begin
              real_value= -29142;
              imag_value=14968;
            end
    1409  : begin
              real_value= -31575;
              imag_value=8737;
            end
    1410  : begin
              real_value= -32691;
              imag_value=2142;
            end
    1411  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    1412  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    1413  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    1414  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    1415  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    1416  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    1417  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    1418  : begin
              real_value= 0;
              imag_value=-32760;
            end
    1419  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    1420  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    1421  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    1422  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    1423  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    1424  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    1425  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    1426  : begin
              real_value= 32691;
              imag_value=2142;
            end
    1427  : begin
              real_value= 31575;
              imag_value=8737;
            end
    1428  : begin
              real_value= 29142;
              imag_value=14968;
            end
    1429  : begin
              real_value= 25494;
              imag_value=20575;
            end
    1430  : begin
              real_value= 20783;
              imag_value=25324;
            end
    1431  : begin
              real_value= 15206;
              imag_value=29017;
            end
    1432  : begin
              real_value= 8995;
              imag_value=31501;
            end
    1433  : begin
              real_value= 2408;
              imag_value=32673;
            end
    1434  : begin
              real_value= -4275;
              imag_value=32481;
            end
    1435  : begin
              real_value= -10783;
              imag_value=30935;
            end
    1436  : begin
              real_value= -16842;
              imag_value=28100;
            end
    1437  : begin
              real_value= -22199;
              imag_value=24092;
            end
    1438  : begin
              real_value= -26630;
              imag_value=19081;
            end
    1439  : begin
              real_value= -29950;
              imag_value=13274;
            end
    1440  : begin
              real_value= -32022;
              imag_value=6915;
            end
    1441  : begin
              real_value= -32759;
              imag_value=267;
            end
    1442  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    1443  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    1444  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    1445  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    1446  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    1447  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    1448  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    1449  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    1450  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    1451  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    1452  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    1453  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    1454  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    1455  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    1456  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    1457  : begin
              real_value= 32515;
              imag_value=4009;
            end
    1458  : begin
              real_value= 31023;
              imag_value=10529;
            end
    1459  : begin
              real_value= 28236;
              imag_value=16611;
            end
    1460  : begin
              real_value= 24274;
              imag_value=22001;
            end
    1461  : begin
              real_value= 19299;
              imag_value=26472;
            end
    1462  : begin
              real_value= 13520;
              imag_value=29841;
            end
    1463  : begin
              real_value= 7177;
              imag_value=31965;
            end
    1464  : begin
              real_value= 535;
              imag_value=32757;
            end
    1465  : begin
              real_value= -6127;
              imag_value=32183;
            end
    1466  : begin
              real_value= -12537;
              imag_value=30267;
            end
    1467  : begin
              real_value= -18423;
              imag_value=27090;
            end
    1468  : begin
              real_value= -23541;
              imag_value=22782;
            end
    1469  : begin
              real_value= -27678;
              imag_value=17525;
            end
    1470  : begin
              real_value= -30661;
              imag_value=11539;
            end
    1471  : begin
              real_value= -32365;
              imag_value=5071;
            end
    1472  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    1473  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    1474  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    1475  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    1476  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    1477  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    1478  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    1479  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    1480  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    1481  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    1482  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    1483  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    1484  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    1485  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    1486  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    1487  : begin
              real_value= 32750;
              imag_value=-802;
            end
    1488  : begin
              real_value= 32231;
              imag_value=5864;
            end
    1489  : begin
              real_value= 30369;
              imag_value=12288;
            end
    1490  : begin
              real_value= 27240;
              imag_value=18200;
            end
    1491  : begin
              real_value= 22974;
              imag_value=23354;
            end
    1492  : begin
              real_value= 17752;
              imag_value=27534;
            end
    1493  : begin
              real_value= 11790;
              imag_value=30565;
            end
    1494  : begin
              real_value= 5336;
              imag_value=32323;
            end
    1495  : begin
              real_value= -1338;
              imag_value=32733;
            end
    1496  : begin
              real_value= -7959;
              imag_value=31779;
            end
    1497  : begin
              real_value= -14248;
              imag_value=29499;
            end
    1498  : begin
              real_value= -19943;
              imag_value=25990;
            end
    1499  : begin
              real_value= -24806;
              imag_value=21399;
            end
    1500  : begin
              real_value= -28636;
              imag_value=15914;
            end
    1501  : begin
              real_value= -31271;
              imag_value=9765;
            end
    1502  : begin
              real_value= -32603;
              imag_value=3210;
            end
    1503  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    1504  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    1505  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    1506  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    1507  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    1508  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    1509  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    1510  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    1511  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    1512  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    1513  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    1514  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    1515  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    1516  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    1517  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    1518  : begin
              real_value= 32743;
              imag_value=1070;
            end
    1519  : begin
              real_value= 31843;
              imag_value=7699;
            end
    1520  : begin
              real_value= 29615;
              imag_value=14006;
            end
    1521  : begin
              real_value= 26152;
              imag_value=19729;
            end
    1522  : begin
              real_value= 21600;
              imag_value=24630;
            end
    1523  : begin
              real_value= 16148;
              imag_value=28506;
            end
    1524  : begin
              real_value= 10021;
              imag_value=31191;
            end
    1525  : begin
              real_value= 3476;
              imag_value=32575;
            end
    1526  : begin
              real_value= -3210;
              imag_value=32603;
            end
    1527  : begin
              real_value= -9765;
              imag_value=31271;
            end
    1528  : begin
              real_value= -15914;
              imag_value=28636;
            end
    1529  : begin
              real_value= -21399;
              imag_value=24806;
            end
    1530  : begin
              real_value= -25990;
              imag_value=19943;
            end
    1531  : begin
              real_value= -29499;
              imag_value=14248;
            end
    1532  : begin
              real_value= -31779;
              imag_value=7959;
            end
    1533  : begin
              real_value= -32733;
              imag_value=1338;
            end
    1534  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    1535  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    1536  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    1537  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    1538  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    1539  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    1540  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    1541  : begin
              real_value= 802;
              imag_value=-32750;
            end
    1542  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    1543  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    1544  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    1545  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    1546  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    1547  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    1548  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    1549  : begin
              real_value= 32629;
              imag_value=2942;
            end
    1550  : begin
              real_value= 31351;
              imag_value=9508;
            end
    1551  : begin
              real_value= 28766;
              imag_value=15678;
            end
    1552  : begin
              real_value= 24981;
              imag_value=21194;
            end
    1553  : begin
              real_value= 20154;
              imag_value=25826;
            end
    1554  : begin
              real_value= 14489;
              imag_value=29382;
            end
    1555  : begin
              real_value= 8219;
              imag_value=31713;
            end
    1556  : begin
              real_value= 1606;
              imag_value=32721;
            end
    1557  : begin
              real_value= -5071;
              imag_value=32365;
            end
    1558  : begin
              real_value= -11539;
              imag_value=30661;
            end
    1559  : begin
              real_value= -17525;
              imag_value=27678;
            end
    1560  : begin
              real_value= -22782;
              imag_value=23541;
            end
    1561  : begin
              real_value= -27090;
              imag_value=18423;
            end
    1562  : begin
              real_value= -30267;
              imag_value=12537;
            end
    1563  : begin
              real_value= -32183;
              imag_value=6127;
            end
    1564  : begin
              real_value= -32757;
              imag_value=-535;
            end
    1565  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    1566  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    1567  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    1568  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    1569  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    1570  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    1571  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    1572  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    1573  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    1574  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    1575  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    1576  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    1577  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    1578  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    1579  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    1580  : begin
              real_value= 32407;
              imag_value=4806;
            end
    1581  : begin
              real_value= 30755;
              imag_value=11289;
            end
    1582  : begin
              real_value= 27820;
              imag_value=17299;
            end
    1583  : begin
              real_value= 23726;
              imag_value=22589;
            end
    1584  : begin
              real_value= 18644;
              imag_value=26938;
            end
    1585  : begin
              real_value= 12784;
              imag_value=30163;
            end
    1586  : begin
              real_value= 6390;
              imag_value=32131;
            end
    1587  : begin
              real_value= -267;
              imag_value=32759;
            end
    1588  : begin
              real_value= -6915;
              imag_value=32022;
            end
    1589  : begin
              real_value= -13274;
              imag_value=29950;
            end
    1590  : begin
              real_value= -19081;
              imag_value=26630;
            end
    1591  : begin
              real_value= -24092;
              imag_value=22199;
            end
    1592  : begin
              real_value= -28100;
              imag_value=16842;
            end
    1593  : begin
              real_value= -30935;
              imag_value=10783;
            end
    1594  : begin
              real_value= -32481;
              imag_value=4275;
            end
    1595  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    1596  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    1597  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    1598  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    1599  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    1600  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    1601  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    1602  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    1603  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    1604  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    1605  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    1606  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    1607  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    1608  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    1609  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    1610  : begin
              real_value= 32760;
              imag_value=0;
            end
    1611  : begin
              real_value= 32077;
              imag_value=6654;
            end
    1612  : begin
              real_value= 30057;
              imag_value=13030;
            end
    1613  : begin
              real_value= 26784;
              imag_value=18863;
            end
    1614  : begin
              real_value= 22395;
              imag_value=23911;
            end
    1615  : begin
              real_value= 17072;
              imag_value=27961;
            end
    1616  : begin
              real_value= 11036;
              imag_value=30846;
            end
    1617  : begin
              real_value= 4540;
              imag_value=32445;
            end
    1618  : begin
              real_value= -2142;
              imag_value=32691;
            end
    1619  : begin
              real_value= -8737;
              imag_value=31575;
            end
    1620  : begin
              real_value= -14968;
              imag_value=29142;
            end
    1621  : begin
              real_value= -20575;
              imag_value=25494;
            end
    1622  : begin
              real_value= -25324;
              imag_value=20783;
            end
    1623  : begin
              real_value= -29017;
              imag_value=15206;
            end
    1624  : begin
              real_value= -31501;
              imag_value=8995;
            end
    1625  : begin
              real_value= -32673;
              imag_value=2408;
            end
    1626  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    1627  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    1628  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    1629  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    1630  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    1631  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    1632  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    1633  : begin
              real_value= -267;
              imag_value=-32759;
            end
    1634  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    1635  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    1636  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    1637  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    1638  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    1639  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    1640  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    1641  : begin
              real_value= 32707;
              imag_value=1874;
            end
    1642  : begin
              real_value= 31645;
              imag_value=8477;
            end
    1643  : begin
              real_value= 29263;
              imag_value=14728;
            end
    1644  : begin
              real_value= 25661;
              imag_value=20365;
            end
    1645  : begin
              real_value= 20988;
              imag_value=25154;
            end
    1646  : begin
              real_value= 15442;
              imag_value=28892;
            end
    1647  : begin
              real_value= 9253;
              imag_value=31426;
            end
    1648  : begin
              real_value= 2676;
              imag_value=32651;
            end
    1649  : begin
              real_value= -4009;
              imag_value=32515;
            end
    1650  : begin
              real_value= -10529;
              imag_value=31023;
            end
    1651  : begin
              real_value= -16611;
              imag_value=28236;
            end
    1652  : begin
              real_value= -22001;
              imag_value=24274;
            end
    1653  : begin
              real_value= -26472;
              imag_value=19299;
            end
    1654  : begin
              real_value= -29841;
              imag_value=13520;
            end
    1655  : begin
              real_value= -31965;
              imag_value=7177;
            end
    1656  : begin
              real_value= -32757;
              imag_value=535;
            end
    1657  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    1658  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    1659  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    1660  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    1661  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    1662  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    1663  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    1664  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    1665  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    1666  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    1667  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    1668  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    1669  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    1670  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    1671  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    1672  : begin
              real_value= 32547;
              imag_value=3742;
            end
    1673  : begin
              real_value= 31107;
              imag_value=10275;
            end
    1674  : begin
              real_value= 28371;
              imag_value=16380;
            end
    1675  : begin
              real_value= 24453;
              imag_value=21801;
            end
    1676  : begin
              real_value= 19515;
              imag_value=26314;
            end
    1677  : begin
              real_value= 13764;
              imag_value=29729;
            end
    1678  : begin
              real_value= 7438;
              imag_value=31905;
            end
    1679  : begin
              real_value= 802;
              imag_value=32750;
            end
    1680  : begin
              real_value= -5864;
              imag_value=32231;
            end
    1681  : begin
              real_value= -12288;
              imag_value=30369;
            end
    1682  : begin
              real_value= -18200;
              imag_value=27240;
            end
    1683  : begin
              real_value= -23354;
              imag_value=22974;
            end
    1684  : begin
              real_value= -27534;
              imag_value=17752;
            end
    1685  : begin
              real_value= -30565;
              imag_value=11790;
            end
    1686  : begin
              real_value= -32323;
              imag_value=5336;
            end
    1687  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    1688  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    1689  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    1690  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    1691  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    1692  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    1693  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    1694  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    1695  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    1696  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    1697  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    1698  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    1699  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    1700  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    1701  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    1702  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    1703  : begin
              real_value= 32278;
              imag_value=5599;
            end
    1704  : begin
              real_value= 30468;
              imag_value=12039;
            end
    1705  : begin
              real_value= 27387;
              imag_value=17977;
            end
    1706  : begin
              real_value= 23165;
              imag_value=23165;
            end
    1707  : begin
              real_value= 17977;
              imag_value=27387;
            end
    1708  : begin
              real_value= 12039;
              imag_value=30468;
            end
    1709  : begin
              real_value= 5599;
              imag_value=32278;
            end
    1710  : begin
              real_value= -1070;
              imag_value=32743;
            end
    1711  : begin
              real_value= -7699;
              imag_value=31843;
            end
    1712  : begin
              real_value= -14006;
              imag_value=29615;
            end
    1713  : begin
              real_value= -19729;
              imag_value=26152;
            end
    1714  : begin
              real_value= -24630;
              imag_value=21600;
            end
    1715  : begin
              real_value= -28506;
              imag_value=16148;
            end
    1716  : begin
              real_value= -31191;
              imag_value=10021;
            end
    1717  : begin
              real_value= -32575;
              imag_value=3476;
            end
    1718  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    1719  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    1720  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    1721  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    1722  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    1723  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    1724  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    1725  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    1726  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    1727  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    1728  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    1729  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    1730  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    1731  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    1732  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    1733  : begin
              real_value= 32750;
              imag_value=802;
            end
    1734  : begin
              real_value= 31905;
              imag_value=7438;
            end
    1735  : begin
              real_value= 29729;
              imag_value=13764;
            end
    1736  : begin
              real_value= 26314;
              imag_value=19515;
            end
    1737  : begin
              real_value= 21801;
              imag_value=24453;
            end
    1738  : begin
              real_value= 16380;
              imag_value=28371;
            end
    1739  : begin
              real_value= 10275;
              imag_value=31107;
            end
    1740  : begin
              real_value= 3742;
              imag_value=32547;
            end
    1741  : begin
              real_value= -2942;
              imag_value=32629;
            end
    1742  : begin
              real_value= -9508;
              imag_value=31351;
            end
    1743  : begin
              real_value= -15678;
              imag_value=28766;
            end
    1744  : begin
              real_value= -21194;
              imag_value=24981;
            end
    1745  : begin
              real_value= -25826;
              imag_value=20154;
            end
    1746  : begin
              real_value= -29382;
              imag_value=14489;
            end
    1747  : begin
              real_value= -31713;
              imag_value=8219;
            end
    1748  : begin
              real_value= -32721;
              imag_value=1606;
            end
    1749  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    1750  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    1751  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    1752  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    1753  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    1754  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    1755  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    1756  : begin
              real_value= 535;
              imag_value=-32757;
            end
    1757  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    1758  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    1759  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    1760  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    1761  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    1762  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    1763  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    1764  : begin
              real_value= 32651;
              imag_value=2676;
            end
    1765  : begin
              real_value= 31426;
              imag_value=9253;
            end
    1766  : begin
              real_value= 28892;
              imag_value=15442;
            end
    1767  : begin
              real_value= 25154;
              imag_value=20988;
            end
    1768  : begin
              real_value= 20365;
              imag_value=25661;
            end
    1769  : begin
              real_value= 14728;
              imag_value=29263;
            end
    1770  : begin
              real_value= 8477;
              imag_value=31645;
            end
    1771  : begin
              real_value= 1874;
              imag_value=32707;
            end
    1772  : begin
              real_value= -4806;
              imag_value=32407;
            end
    1773  : begin
              real_value= -11289;
              imag_value=30755;
            end
    1774  : begin
              real_value= -17299;
              imag_value=27820;
            end
    1775  : begin
              real_value= -22589;
              imag_value=23726;
            end
    1776  : begin
              real_value= -26938;
              imag_value=18644;
            end
    1777  : begin
              real_value= -30163;
              imag_value=12784;
            end
    1778  : begin
              real_value= -32131;
              imag_value=6390;
            end
    1779  : begin
              real_value= -32759;
              imag_value=-267;
            end
    1780  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    1781  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    1782  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    1783  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    1784  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    1785  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    1786  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    1787  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    1788  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    1789  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    1790  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    1791  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    1792  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    1793  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    1794  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    1795  : begin
              real_value= 32445;
              imag_value=4540;
            end
    1796  : begin
              real_value= 30846;
              imag_value=11036;
            end
    1797  : begin
              real_value= 27961;
              imag_value=17072;
            end
    1798  : begin
              real_value= 23911;
              imag_value=22395;
            end
    1799  : begin
              real_value= 18863;
              imag_value=26784;
            end
    1800  : begin
              real_value= 13030;
              imag_value=30057;
            end
    1801  : begin
              real_value= 6654;
              imag_value=32077;
            end
    1802  : begin
              real_value= 0;
              imag_value=32760;
            end
    1803  : begin
              real_value= -6654;
              imag_value=32077;
            end
    1804  : begin
              real_value= -13030;
              imag_value=30057;
            end
    1805  : begin
              real_value= -18863;
              imag_value=26784;
            end
    1806  : begin
              real_value= -23911;
              imag_value=22395;
            end
    1807  : begin
              real_value= -27961;
              imag_value=17072;
            end
    1808  : begin
              real_value= -30846;
              imag_value=11036;
            end
    1809  : begin
              real_value= -32445;
              imag_value=4540;
            end
    1810  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    1811  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    1812  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    1813  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    1814  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    1815  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    1816  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    1817  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    1818  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    1819  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    1820  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    1821  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    1822  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    1823  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    1824  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    1825  : begin
              real_value= 32759;
              imag_value=-267;
            end
    1826  : begin
              real_value= 32131;
              imag_value=6390;
            end
    1827  : begin
              real_value= 30163;
              imag_value=12784;
            end
    1828  : begin
              real_value= 26938;
              imag_value=18644;
            end
    1829  : begin
              real_value= 22589;
              imag_value=23726;
            end
    1830  : begin
              real_value= 17299;
              imag_value=27820;
            end
    1831  : begin
              real_value= 11289;
              imag_value=30755;
            end
    1832  : begin
              real_value= 4806;
              imag_value=32407;
            end
    1833  : begin
              real_value= -1874;
              imag_value=32707;
            end
    1834  : begin
              real_value= -8477;
              imag_value=31645;
            end
    1835  : begin
              real_value= -14728;
              imag_value=29263;
            end
    1836  : begin
              real_value= -20365;
              imag_value=25661;
            end
    1837  : begin
              real_value= -25154;
              imag_value=20988;
            end
    1838  : begin
              real_value= -28892;
              imag_value=15442;
            end
    1839  : begin
              real_value= -31426;
              imag_value=9253;
            end
    1840  : begin
              real_value= -32651;
              imag_value=2676;
            end
    1841  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    1842  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    1843  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    1844  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    1845  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    1846  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    1847  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    1848  : begin
              real_value= -535;
              imag_value=-32757;
            end
    1849  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    1850  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    1851  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    1852  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    1853  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    1854  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    1855  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    1856  : begin
              real_value= 32721;
              imag_value=1606;
            end
    1857  : begin
              real_value= 31713;
              imag_value=8219;
            end
    1858  : begin
              real_value= 29382;
              imag_value=14489;
            end
    1859  : begin
              real_value= 25826;
              imag_value=20154;
            end
    1860  : begin
              real_value= 21194;
              imag_value=24981;
            end
    1861  : begin
              real_value= 15678;
              imag_value=28766;
            end
    1862  : begin
              real_value= 9508;
              imag_value=31351;
            end
    1863  : begin
              real_value= 2942;
              imag_value=32629;
            end
    1864  : begin
              real_value= -3742;
              imag_value=32547;
            end
    1865  : begin
              real_value= -10275;
              imag_value=31107;
            end
    1866  : begin
              real_value= -16380;
              imag_value=28371;
            end
    1867  : begin
              real_value= -21801;
              imag_value=24453;
            end
    1868  : begin
              real_value= -26314;
              imag_value=19515;
            end
    1869  : begin
              real_value= -29729;
              imag_value=13764;
            end
    1870  : begin
              real_value= -31905;
              imag_value=7438;
            end
    1871  : begin
              real_value= -32750;
              imag_value=802;
            end
    1872  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    1873  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    1874  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    1875  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    1876  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    1877  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    1878  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    1879  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    1880  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    1881  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    1882  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    1883  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    1884  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    1885  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    1886  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    1887  : begin
              real_value= 32575;
              imag_value=3476;
            end
    1888  : begin
              real_value= 31191;
              imag_value=10021;
            end
    1889  : begin
              real_value= 28506;
              imag_value=16148;
            end
    1890  : begin
              real_value= 24630;
              imag_value=21600;
            end
    1891  : begin
              real_value= 19729;
              imag_value=26152;
            end
    1892  : begin
              real_value= 14006;
              imag_value=29615;
            end
    1893  : begin
              real_value= 7699;
              imag_value=31843;
            end
    1894  : begin
              real_value= 1070;
              imag_value=32743;
            end
    1895  : begin
              real_value= -5599;
              imag_value=32278;
            end
    1896  : begin
              real_value= -12039;
              imag_value=30468;
            end
    1897  : begin
              real_value= -17977;
              imag_value=27387;
            end
    1898  : begin
              real_value= -23165;
              imag_value=23165;
            end
    1899  : begin
              real_value= -27387;
              imag_value=17977;
            end
    1900  : begin
              real_value= -30468;
              imag_value=12039;
            end
    1901  : begin
              real_value= -32278;
              imag_value=5599;
            end
    1902  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    1903  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    1904  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    1905  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    1906  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    1907  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    1908  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    1909  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    1910  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    1911  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    1912  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    1913  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    1914  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    1915  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    1916  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    1917  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    1918  : begin
              real_value= 32323;
              imag_value=5336;
            end
    1919  : begin
              real_value= 30565;
              imag_value=11790;
            end
    1920  : begin
              real_value= 27534;
              imag_value=17752;
            end
    1921  : begin
              real_value= 23354;
              imag_value=22974;
            end
    1922  : begin
              real_value= 18200;
              imag_value=27240;
            end
    1923  : begin
              real_value= 12288;
              imag_value=30369;
            end
    1924  : begin
              real_value= 5864;
              imag_value=32231;
            end
    1925  : begin
              real_value= -802;
              imag_value=32750;
            end
    1926  : begin
              real_value= -7438;
              imag_value=31905;
            end
    1927  : begin
              real_value= -13764;
              imag_value=29729;
            end
    1928  : begin
              real_value= -19515;
              imag_value=26314;
            end
    1929  : begin
              real_value= -24453;
              imag_value=21801;
            end
    1930  : begin
              real_value= -28371;
              imag_value=16380;
            end
    1931  : begin
              real_value= -31107;
              imag_value=10275;
            end
    1932  : begin
              real_value= -32547;
              imag_value=3742;
            end
    1933  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    1934  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    1935  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    1936  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    1937  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    1938  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    1939  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    1940  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    1941  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    1942  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    1943  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    1944  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    1945  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    1946  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    1947  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    1948  : begin
              real_value= 32757;
              imag_value=535;
            end
    1949  : begin
              real_value= 31965;
              imag_value=7177;
            end
    1950  : begin
              real_value= 29841;
              imag_value=13520;
            end
    1951  : begin
              real_value= 26472;
              imag_value=19299;
            end
    1952  : begin
              real_value= 22001;
              imag_value=24274;
            end
    1953  : begin
              real_value= 16611;
              imag_value=28236;
            end
    1954  : begin
              real_value= 10529;
              imag_value=31023;
            end
    1955  : begin
              real_value= 4009;
              imag_value=32515;
            end
    1956  : begin
              real_value= -2676;
              imag_value=32651;
            end
    1957  : begin
              real_value= -9253;
              imag_value=31426;
            end
    1958  : begin
              real_value= -15442;
              imag_value=28892;
            end
    1959  : begin
              real_value= -20988;
              imag_value=25154;
            end
    1960  : begin
              real_value= -25661;
              imag_value=20365;
            end
    1961  : begin
              real_value= -29263;
              imag_value=14728;
            end
    1962  : begin
              real_value= -31645;
              imag_value=8477;
            end
    1963  : begin
              real_value= -32707;
              imag_value=1874;
            end
    1964  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    1965  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    1966  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    1967  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    1968  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    1969  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    1970  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    1971  : begin
              real_value= 267;
              imag_value=-32759;
            end
    1972  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    1973  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    1974  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    1975  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    1976  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    1977  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    1978  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    1979  : begin
              real_value= 32673;
              imag_value=2408;
            end
    1980  : begin
              real_value= 31501;
              imag_value=8995;
            end
    1981  : begin
              real_value= 29017;
              imag_value=15206;
            end
    1982  : begin
              real_value= 25324;
              imag_value=20783;
            end
    1983  : begin
              real_value= 20575;
              imag_value=25494;
            end
    1984  : begin
              real_value= 14968;
              imag_value=29142;
            end
    1985  : begin
              real_value= 8737;
              imag_value=31575;
            end
    1986  : begin
              real_value= 2142;
              imag_value=32691;
            end
    1987  : begin
              real_value= -4540;
              imag_value=32445;
            end
    1988  : begin
              real_value= -11036;
              imag_value=30846;
            end
    1989  : begin
              real_value= -17072;
              imag_value=27961;
            end
    1990  : begin
              real_value= -22395;
              imag_value=23911;
            end
    1991  : begin
              real_value= -26784;
              imag_value=18863;
            end
    1992  : begin
              real_value= -30057;
              imag_value=13030;
            end
    1993  : begin
              real_value= -32077;
              imag_value=6654;
            end
    1994  : begin
              real_value= -32760;
              imag_value=0;
            end
    1995  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    1996  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    1997  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    1998  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    1999  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    2000  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    2001  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    2002  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    2003  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    2004  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    2005  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    2006  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    2007  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    2008  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    2009  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    2010  : begin
              real_value= 32481;
              imag_value=4275;
            end
    2011  : begin
              real_value= 30935;
              imag_value=10783;
            end
    2012  : begin
              real_value= 28100;
              imag_value=16842;
            end
    2013  : begin
              real_value= 24092;
              imag_value=22199;
            end
    2014  : begin
              real_value= 19081;
              imag_value=26630;
            end
    2015  : begin
              real_value= 13274;
              imag_value=29950;
            end
    2016  : begin
              real_value= 6915;
              imag_value=32022;
            end
    2017  : begin
              real_value= 267;
              imag_value=32759;
            end
    2018  : begin
              real_value= -6390;
              imag_value=32131;
            end
    2019  : begin
              real_value= -12784;
              imag_value=30163;
            end
    2020  : begin
              real_value= -18644;
              imag_value=26938;
            end
    2021  : begin
              real_value= -23726;
              imag_value=22589;
            end
    2022  : begin
              real_value= -27820;
              imag_value=17299;
            end
    2023  : begin
              real_value= -30755;
              imag_value=11289;
            end
    2024  : begin
              real_value= -32407;
              imag_value=4806;
            end
    2025  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    2026  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    2027  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    2028  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    2029  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    2030  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    2031  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    2032  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    2033  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    2034  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    2035  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    2036  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    2037  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    2038  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    2039  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    2040  : begin
              real_value= 32757;
              imag_value=-535;
            end
    2041  : begin
              real_value= 32183;
              imag_value=6127;
            end
    2042  : begin
              real_value= 30267;
              imag_value=12537;
            end
    2043  : begin
              real_value= 27090;
              imag_value=18423;
            end
    2044  : begin
              real_value= 22782;
              imag_value=23541;
            end
    2045  : begin
              real_value= 17525;
              imag_value=27678;
            end
    2046  : begin
              real_value= 11539;
              imag_value=30661;
            end
    2047  : begin
              real_value= 5071;
              imag_value=32365;
            end
    2048  : begin
              real_value= -1606;
              imag_value=32721;
            end
    2049  : begin
              real_value= -8219;
              imag_value=31713;
            end
    2050  : begin
              real_value= -14489;
              imag_value=29382;
            end
    2051  : begin
              real_value= -20154;
              imag_value=25826;
            end
    2052  : begin
              real_value= -24981;
              imag_value=21194;
            end
    2053  : begin
              real_value= -28766;
              imag_value=15678;
            end
    2054  : begin
              real_value= -31351;
              imag_value=9508;
            end
    2055  : begin
              real_value= -32629;
              imag_value=2942;
            end
    2056  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    2057  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    2058  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    2059  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    2060  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    2061  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    2062  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    2063  : begin
              real_value= -802;
              imag_value=-32750;
            end
    2064  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    2065  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    2066  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    2067  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    2068  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    2069  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    2070  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    2071  : begin
              real_value= 32733;
              imag_value=1338;
            end
    2072  : begin
              real_value= 31779;
              imag_value=7959;
            end
    2073  : begin
              real_value= 29499;
              imag_value=14248;
            end
    2074  : begin
              real_value= 25990;
              imag_value=19943;
            end
    2075  : begin
              real_value= 21399;
              imag_value=24806;
            end
    2076  : begin
              real_value= 15914;
              imag_value=28636;
            end
    2077  : begin
              real_value= 9765;
              imag_value=31271;
            end
    2078  : begin
              real_value= 3210;
              imag_value=32603;
            end
    2079  : begin
              real_value= -3476;
              imag_value=32575;
            end
    2080  : begin
              real_value= -10021;
              imag_value=31191;
            end
    2081  : begin
              real_value= -16148;
              imag_value=28506;
            end
    2082  : begin
              real_value= -21600;
              imag_value=24630;
            end
    2083  : begin
              real_value= -26152;
              imag_value=19729;
            end
    2084  : begin
              real_value= -29615;
              imag_value=14006;
            end
    2085  : begin
              real_value= -31843;
              imag_value=7699;
            end
    2086  : begin
              real_value= -32743;
              imag_value=1070;
            end
    2087  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    2088  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    2089  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    2090  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    2091  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    2092  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    2093  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    2094  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    2095  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    2096  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    2097  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    2098  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    2099  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    2100  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    2101  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    2102  : begin
              real_value= 32603;
              imag_value=3210;
            end
    2103  : begin
              real_value= 31271;
              imag_value=9765;
            end
    2104  : begin
              real_value= 28636;
              imag_value=15914;
            end
    2105  : begin
              real_value= 24806;
              imag_value=21399;
            end
    2106  : begin
              real_value= 19943;
              imag_value=25990;
            end
    2107  : begin
              real_value= 14248;
              imag_value=29499;
            end
    2108  : begin
              real_value= 7959;
              imag_value=31779;
            end
    2109  : begin
              real_value= 1338;
              imag_value=32733;
            end
    2110  : begin
              real_value= -5336;
              imag_value=32323;
            end
    2111  : begin
              real_value= -11790;
              imag_value=30565;
            end
    2112  : begin
              real_value= -17752;
              imag_value=27534;
            end
    2113  : begin
              real_value= -22974;
              imag_value=23354;
            end
    2114  : begin
              real_value= -27240;
              imag_value=18200;
            end
    2115  : begin
              real_value= -30369;
              imag_value=12288;
            end
    2116  : begin
              real_value= -32231;
              imag_value=5864;
            end
    2117  : begin
              real_value= -32750;
              imag_value=-802;
            end
    2118  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    2119  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    2120  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    2121  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    2122  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    2123  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    2124  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    2125  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    2126  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    2127  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    2128  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    2129  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    2130  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    2131  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    2132  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    2133  : begin
              real_value= 32365;
              imag_value=5071;
            end
    2134  : begin
              real_value= 30661;
              imag_value=11539;
            end
    2135  : begin
              real_value= 27678;
              imag_value=17525;
            end
    2136  : begin
              real_value= 23541;
              imag_value=22782;
            end
    2137  : begin
              real_value= 18423;
              imag_value=27090;
            end
    2138  : begin
              real_value= 12537;
              imag_value=30267;
            end
    2139  : begin
              real_value= 6127;
              imag_value=32183;
            end
    2140  : begin
              real_value= -535;
              imag_value=32757;
            end
    2141  : begin
              real_value= -7177;
              imag_value=31965;
            end
    2142  : begin
              real_value= -13520;
              imag_value=29841;
            end
    2143  : begin
              real_value= -19299;
              imag_value=26472;
            end
    2144  : begin
              real_value= -24274;
              imag_value=22001;
            end
    2145  : begin
              real_value= -28236;
              imag_value=16611;
            end
    2146  : begin
              real_value= -31023;
              imag_value=10529;
            end
    2147  : begin
              real_value= -32515;
              imag_value=4009;
            end
    2148  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    2149  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    2150  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    2151  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    2152  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    2153  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    2154  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    2155  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    2156  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    2157  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    2158  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    2159  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    2160  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    2161  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    2162  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    2163  : begin
              real_value= 32759;
              imag_value=267;
            end
    2164  : begin
              real_value= 32022;
              imag_value=6915;
            end
    2165  : begin
              real_value= 29950;
              imag_value=13274;
            end
    2166  : begin
              real_value= 26630;
              imag_value=19081;
            end
    2167  : begin
              real_value= 22199;
              imag_value=24092;
            end
    2168  : begin
              real_value= 16842;
              imag_value=28100;
            end
    2169  : begin
              real_value= 10783;
              imag_value=30935;
            end
    2170  : begin
              real_value= 4275;
              imag_value=32481;
            end
    2171  : begin
              real_value= -2408;
              imag_value=32673;
            end
    2172  : begin
              real_value= -8995;
              imag_value=31501;
            end
    2173  : begin
              real_value= -15206;
              imag_value=29017;
            end
    2174  : begin
              real_value= -20783;
              imag_value=25324;
            end
    2175  : begin
              real_value= -25494;
              imag_value=20575;
            end
    2176  : begin
              real_value= -29142;
              imag_value=14968;
            end
    2177  : begin
              real_value= -31575;
              imag_value=8737;
            end
    2178  : begin
              real_value= -32691;
              imag_value=2142;
            end
    2179  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    2180  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    2181  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    2182  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    2183  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    2184  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    2185  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    2186  : begin
              real_value= 0;
              imag_value=-32760;
            end
    2187  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    2188  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    2189  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    2190  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    2191  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    2192  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    2193  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    2194  : begin
              real_value= 32691;
              imag_value=2142;
            end
    2195  : begin
              real_value= 31575;
              imag_value=8737;
            end
    2196  : begin
              real_value= 29142;
              imag_value=14968;
            end
    2197  : begin
              real_value= 25494;
              imag_value=20575;
            end
    2198  : begin
              real_value= 20783;
              imag_value=25324;
            end
    2199  : begin
              real_value= 15206;
              imag_value=29017;
            end
    2200  : begin
              real_value= 8995;
              imag_value=31501;
            end
    2201  : begin
              real_value= 2408;
              imag_value=32673;
            end
    2202  : begin
              real_value= -4275;
              imag_value=32481;
            end
    2203  : begin
              real_value= -10783;
              imag_value=30935;
            end
    2204  : begin
              real_value= -16842;
              imag_value=28100;
            end
    2205  : begin
              real_value= -22199;
              imag_value=24092;
            end
    2206  : begin
              real_value= -26630;
              imag_value=19081;
            end
    2207  : begin
              real_value= -29950;
              imag_value=13274;
            end
    2208  : begin
              real_value= -32022;
              imag_value=6915;
            end
    2209  : begin
              real_value= -32759;
              imag_value=267;
            end
    2210  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    2211  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    2212  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    2213  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    2214  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    2215  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    2216  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    2217  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    2218  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    2219  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    2220  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    2221  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    2222  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    2223  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    2224  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    2225  : begin
              real_value= 32515;
              imag_value=4009;
            end
    2226  : begin
              real_value= 31023;
              imag_value=10529;
            end
    2227  : begin
              real_value= 28236;
              imag_value=16611;
            end
    2228  : begin
              real_value= 24274;
              imag_value=22001;
            end
    2229  : begin
              real_value= 19299;
              imag_value=26472;
            end
    2230  : begin
              real_value= 13520;
              imag_value=29841;
            end
    2231  : begin
              real_value= 7177;
              imag_value=31965;
            end
    2232  : begin
              real_value= 535;
              imag_value=32757;
            end
    2233  : begin
              real_value= -6127;
              imag_value=32183;
            end
    2234  : begin
              real_value= -12537;
              imag_value=30267;
            end
    2235  : begin
              real_value= -18423;
              imag_value=27090;
            end
    2236  : begin
              real_value= -23541;
              imag_value=22782;
            end
    2237  : begin
              real_value= -27678;
              imag_value=17525;
            end
    2238  : begin
              real_value= -30661;
              imag_value=11539;
            end
    2239  : begin
              real_value= -32365;
              imag_value=5071;
            end
    2240  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    2241  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    2242  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    2243  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    2244  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    2245  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    2246  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    2247  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    2248  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    2249  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    2250  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    2251  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    2252  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    2253  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    2254  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    2255  : begin
              real_value= 32750;
              imag_value=-802;
            end
    2256  : begin
              real_value= 32231;
              imag_value=5864;
            end
    2257  : begin
              real_value= 30369;
              imag_value=12288;
            end
    2258  : begin
              real_value= 27240;
              imag_value=18200;
            end
    2259  : begin
              real_value= 22974;
              imag_value=23354;
            end
    2260  : begin
              real_value= 17752;
              imag_value=27534;
            end
    2261  : begin
              real_value= 11790;
              imag_value=30565;
            end
    2262  : begin
              real_value= 5336;
              imag_value=32323;
            end
    2263  : begin
              real_value= -1338;
              imag_value=32733;
            end
    2264  : begin
              real_value= -7959;
              imag_value=31779;
            end
    2265  : begin
              real_value= -14248;
              imag_value=29499;
            end
    2266  : begin
              real_value= -19943;
              imag_value=25990;
            end
    2267  : begin
              real_value= -24806;
              imag_value=21399;
            end
    2268  : begin
              real_value= -28636;
              imag_value=15914;
            end
    2269  : begin
              real_value= -31271;
              imag_value=9765;
            end
    2270  : begin
              real_value= -32603;
              imag_value=3210;
            end
    2271  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    2272  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    2273  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    2274  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    2275  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    2276  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    2277  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    2278  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    2279  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    2280  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    2281  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    2282  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    2283  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    2284  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    2285  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    2286  : begin
              real_value= 32743;
              imag_value=1070;
            end
    2287  : begin
              real_value= 31843;
              imag_value=7699;
            end
    2288  : begin
              real_value= 29615;
              imag_value=14006;
            end
    2289  : begin
              real_value= 26152;
              imag_value=19729;
            end
    2290  : begin
              real_value= 21600;
              imag_value=24630;
            end
    2291  : begin
              real_value= 16148;
              imag_value=28506;
            end
    2292  : begin
              real_value= 10021;
              imag_value=31191;
            end
    2293  : begin
              real_value= 3476;
              imag_value=32575;
            end
    2294  : begin
              real_value= -3210;
              imag_value=32603;
            end
    2295  : begin
              real_value= -9765;
              imag_value=31271;
            end
    2296  : begin
              real_value= -15914;
              imag_value=28636;
            end
    2297  : begin
              real_value= -21399;
              imag_value=24806;
            end
    2298  : begin
              real_value= -25990;
              imag_value=19943;
            end
    2299  : begin
              real_value= -29499;
              imag_value=14248;
            end
    2300  : begin
              real_value= -31779;
              imag_value=7959;
            end
    2301  : begin
              real_value= -32733;
              imag_value=1338;
            end
    2302  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    2303  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    2304  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    2305  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    2306  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    2307  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    2308  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    2309  : begin
              real_value= 802;
              imag_value=-32750;
            end
    2310  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    2311  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    2312  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    2313  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    2314  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    2315  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    2316  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    2317  : begin
              real_value= 32629;
              imag_value=2942;
            end
    2318  : begin
              real_value= 31351;
              imag_value=9508;
            end
    2319  : begin
              real_value= 28766;
              imag_value=15678;
            end
    2320  : begin
              real_value= 24981;
              imag_value=21194;
            end
    2321  : begin
              real_value= 20154;
              imag_value=25826;
            end
    2322  : begin
              real_value= 14489;
              imag_value=29382;
            end
    2323  : begin
              real_value= 8219;
              imag_value=31713;
            end
    2324  : begin
              real_value= 1606;
              imag_value=32721;
            end
    2325  : begin
              real_value= -5071;
              imag_value=32365;
            end
    2326  : begin
              real_value= -11539;
              imag_value=30661;
            end
    2327  : begin
              real_value= -17525;
              imag_value=27678;
            end
    2328  : begin
              real_value= -22782;
              imag_value=23541;
            end
    2329  : begin
              real_value= -27090;
              imag_value=18423;
            end
    2330  : begin
              real_value= -30267;
              imag_value=12537;
            end
    2331  : begin
              real_value= -32183;
              imag_value=6127;
            end
    2332  : begin
              real_value= -32757;
              imag_value=-535;
            end
    2333  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    2334  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    2335  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    2336  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    2337  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    2338  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    2339  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    2340  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    2341  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    2342  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    2343  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    2344  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    2345  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    2346  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    2347  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    2348  : begin
              real_value= 32407;
              imag_value=4806;
            end
    2349  : begin
              real_value= 30755;
              imag_value=11289;
            end
    2350  : begin
              real_value= 27820;
              imag_value=17299;
            end
    2351  : begin
              real_value= 23726;
              imag_value=22589;
            end
    2352  : begin
              real_value= 18644;
              imag_value=26938;
            end
    2353  : begin
              real_value= 12784;
              imag_value=30163;
            end
    2354  : begin
              real_value= 6390;
              imag_value=32131;
            end
    2355  : begin
              real_value= -267;
              imag_value=32759;
            end
    2356  : begin
              real_value= -6915;
              imag_value=32022;
            end
    2357  : begin
              real_value= -13274;
              imag_value=29950;
            end
    2358  : begin
              real_value= -19081;
              imag_value=26630;
            end
    2359  : begin
              real_value= -24092;
              imag_value=22199;
            end
    2360  : begin
              real_value= -28100;
              imag_value=16842;
            end
    2361  : begin
              real_value= -30935;
              imag_value=10783;
            end
    2362  : begin
              real_value= -32481;
              imag_value=4275;
            end
    2363  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    2364  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    2365  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    2366  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    2367  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    2368  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    2369  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    2370  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    2371  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    2372  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    2373  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    2374  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    2375  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    2376  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    2377  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    2378  : begin
              real_value= 32760;
              imag_value=0;
            end
    2379  : begin
              real_value= 32077;
              imag_value=6654;
            end
    2380  : begin
              real_value= 30057;
              imag_value=13030;
            end
    2381  : begin
              real_value= 26784;
              imag_value=18863;
            end
    2382  : begin
              real_value= 22395;
              imag_value=23911;
            end
    2383  : begin
              real_value= 17072;
              imag_value=27961;
            end
    2384  : begin
              real_value= 11036;
              imag_value=30846;
            end
    2385  : begin
              real_value= 4540;
              imag_value=32445;
            end
    2386  : begin
              real_value= -2142;
              imag_value=32691;
            end
    2387  : begin
              real_value= -8737;
              imag_value=31575;
            end
    2388  : begin
              real_value= -14968;
              imag_value=29142;
            end
    2389  : begin
              real_value= -20575;
              imag_value=25494;
            end
    2390  : begin
              real_value= -25324;
              imag_value=20783;
            end
    2391  : begin
              real_value= -29017;
              imag_value=15206;
            end
    2392  : begin
              real_value= -31501;
              imag_value=8995;
            end
    2393  : begin
              real_value= -32673;
              imag_value=2408;
            end
    2394  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    2395  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    2396  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    2397  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    2398  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    2399  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    2400  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    2401  : begin
              real_value= -267;
              imag_value=-32759;
            end
    2402  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    2403  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    2404  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    2405  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    2406  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    2407  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    2408  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    2409  : begin
              real_value= 32707;
              imag_value=1874;
            end
    2410  : begin
              real_value= 31645;
              imag_value=8477;
            end
    2411  : begin
              real_value= 29263;
              imag_value=14728;
            end
    2412  : begin
              real_value= 25661;
              imag_value=20365;
            end
    2413  : begin
              real_value= 20988;
              imag_value=25154;
            end
    2414  : begin
              real_value= 15442;
              imag_value=28892;
            end
    2415  : begin
              real_value= 9253;
              imag_value=31426;
            end
    2416  : begin
              real_value= 2676;
              imag_value=32651;
            end
    2417  : begin
              real_value= -4009;
              imag_value=32515;
            end
    2418  : begin
              real_value= -10529;
              imag_value=31023;
            end
    2419  : begin
              real_value= -16611;
              imag_value=28236;
            end
    2420  : begin
              real_value= -22001;
              imag_value=24274;
            end
    2421  : begin
              real_value= -26472;
              imag_value=19299;
            end
    2422  : begin
              real_value= -29841;
              imag_value=13520;
            end
    2423  : begin
              real_value= -31965;
              imag_value=7177;
            end
    2424  : begin
              real_value= -32757;
              imag_value=535;
            end
    2425  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    2426  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    2427  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    2428  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    2429  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    2430  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    2431  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    2432  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    2433  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    2434  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    2435  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    2436  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    2437  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    2438  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    2439  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    2440  : begin
              real_value= 32547;
              imag_value=3742;
            end
    2441  : begin
              real_value= 31107;
              imag_value=10275;
            end
    2442  : begin
              real_value= 28371;
              imag_value=16380;
            end
    2443  : begin
              real_value= 24453;
              imag_value=21801;
            end
    2444  : begin
              real_value= 19515;
              imag_value=26314;
            end
    2445  : begin
              real_value= 13764;
              imag_value=29729;
            end
    2446  : begin
              real_value= 7438;
              imag_value=31905;
            end
    2447  : begin
              real_value= 802;
              imag_value=32750;
            end
    2448  : begin
              real_value= -5864;
              imag_value=32231;
            end
    2449  : begin
              real_value= -12288;
              imag_value=30369;
            end
    2450  : begin
              real_value= -18200;
              imag_value=27240;
            end
    2451  : begin
              real_value= -23354;
              imag_value=22974;
            end
    2452  : begin
              real_value= -27534;
              imag_value=17752;
            end
    2453  : begin
              real_value= -30565;
              imag_value=11790;
            end
    2454  : begin
              real_value= -32323;
              imag_value=5336;
            end
    2455  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    2456  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    2457  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    2458  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    2459  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    2460  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    2461  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    2462  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    2463  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    2464  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    2465  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    2466  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    2467  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    2468  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    2469  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    2470  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    2471  : begin
              real_value= 32278;
              imag_value=5599;
            end
    2472  : begin
              real_value= 30468;
              imag_value=12039;
            end
    2473  : begin
              real_value= 27387;
              imag_value=17977;
            end
    2474  : begin
              real_value= 23165;
              imag_value=23165;
            end
    2475  : begin
              real_value= 17977;
              imag_value=27387;
            end
    2476  : begin
              real_value= 12039;
              imag_value=30468;
            end
    2477  : begin
              real_value= 5599;
              imag_value=32278;
            end
    2478  : begin
              real_value= -1070;
              imag_value=32743;
            end
    2479  : begin
              real_value= -7699;
              imag_value=31843;
            end
    2480  : begin
              real_value= -14006;
              imag_value=29615;
            end
    2481  : begin
              real_value= -19729;
              imag_value=26152;
            end
    2482  : begin
              real_value= -24630;
              imag_value=21600;
            end
    2483  : begin
              real_value= -28506;
              imag_value=16148;
            end
    2484  : begin
              real_value= -31191;
              imag_value=10021;
            end
    2485  : begin
              real_value= -32575;
              imag_value=3476;
            end
    2486  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    2487  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    2488  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    2489  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    2490  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    2491  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    2492  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    2493  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    2494  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    2495  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    2496  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    2497  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    2498  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    2499  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    2500  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    2501  : begin
              real_value= 32750;
              imag_value=802;
            end
    2502  : begin
              real_value= 31905;
              imag_value=7438;
            end
    2503  : begin
              real_value= 29729;
              imag_value=13764;
            end
    2504  : begin
              real_value= 26314;
              imag_value=19515;
            end
    2505  : begin
              real_value= 21801;
              imag_value=24453;
            end
    2506  : begin
              real_value= 16380;
              imag_value=28371;
            end
    2507  : begin
              real_value= 10275;
              imag_value=31107;
            end
    2508  : begin
              real_value= 3742;
              imag_value=32547;
            end
    2509  : begin
              real_value= -2942;
              imag_value=32629;
            end
    2510  : begin
              real_value= -9508;
              imag_value=31351;
            end
    2511  : begin
              real_value= -15678;
              imag_value=28766;
            end
    2512  : begin
              real_value= -21194;
              imag_value=24981;
            end
    2513  : begin
              real_value= -25826;
              imag_value=20154;
            end
    2514  : begin
              real_value= -29382;
              imag_value=14489;
            end
    2515  : begin
              real_value= -31713;
              imag_value=8219;
            end
    2516  : begin
              real_value= -32721;
              imag_value=1606;
            end
    2517  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    2518  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    2519  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    2520  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    2521  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    2522  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    2523  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    2524  : begin
              real_value= 535;
              imag_value=-32757;
            end
    2525  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    2526  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    2527  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    2528  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    2529  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    2530  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    2531  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    2532  : begin
              real_value= 32651;
              imag_value=2676;
            end
    2533  : begin
              real_value= 31426;
              imag_value=9253;
            end
    2534  : begin
              real_value= 28892;
              imag_value=15442;
            end
    2535  : begin
              real_value= 25154;
              imag_value=20988;
            end
    2536  : begin
              real_value= 20365;
              imag_value=25661;
            end
    2537  : begin
              real_value= 14728;
              imag_value=29263;
            end
    2538  : begin
              real_value= 8477;
              imag_value=31645;
            end
    2539  : begin
              real_value= 1874;
              imag_value=32707;
            end
    2540  : begin
              real_value= -4806;
              imag_value=32407;
            end
    2541  : begin
              real_value= -11289;
              imag_value=30755;
            end
    2542  : begin
              real_value= -17299;
              imag_value=27820;
            end
    2543  : begin
              real_value= -22589;
              imag_value=23726;
            end
    2544  : begin
              real_value= -26938;
              imag_value=18644;
            end
    2545  : begin
              real_value= -30163;
              imag_value=12784;
            end
    2546  : begin
              real_value= -32131;
              imag_value=6390;
            end
    2547  : begin
              real_value= -32759;
              imag_value=-267;
            end
    2548  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    2549  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    2550  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    2551  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    2552  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    2553  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    2554  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    2555  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    2556  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    2557  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    2558  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    2559  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    2560  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    2561  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    2562  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    2563  : begin
              real_value= 32445;
              imag_value=4540;
            end
    2564  : begin
              real_value= 30846;
              imag_value=11036;
            end
    2565  : begin
              real_value= 27961;
              imag_value=17072;
            end
    2566  : begin
              real_value= 23911;
              imag_value=22395;
            end
    2567  : begin
              real_value= 18863;
              imag_value=26784;
            end
    2568  : begin
              real_value= 13030;
              imag_value=30057;
            end
    2569  : begin
              real_value= 6654;
              imag_value=32077;
            end
    2570  : begin
              real_value= 0;
              imag_value=32760;
            end
    2571  : begin
              real_value= -6654;
              imag_value=32077;
            end
    2572  : begin
              real_value= -13030;
              imag_value=30057;
            end
    2573  : begin
              real_value= -18863;
              imag_value=26784;
            end
    2574  : begin
              real_value= -23911;
              imag_value=22395;
            end
    2575  : begin
              real_value= -27961;
              imag_value=17072;
            end
    2576  : begin
              real_value= -30846;
              imag_value=11036;
            end
    2577  : begin
              real_value= -32445;
              imag_value=4540;
            end
    2578  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    2579  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    2580  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    2581  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    2582  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    2583  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    2584  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    2585  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    2586  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    2587  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    2588  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    2589  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    2590  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    2591  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    2592  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    2593  : begin
              real_value= 32759;
              imag_value=-267;
            end
    2594  : begin
              real_value= 32131;
              imag_value=6390;
            end
    2595  : begin
              real_value= 30163;
              imag_value=12784;
            end
    2596  : begin
              real_value= 26938;
              imag_value=18644;
            end
    2597  : begin
              real_value= 22589;
              imag_value=23726;
            end
    2598  : begin
              real_value= 17299;
              imag_value=27820;
            end
    2599  : begin
              real_value= 11289;
              imag_value=30755;
            end
    2600  : begin
              real_value= 4806;
              imag_value=32407;
            end
    2601  : begin
              real_value= -1874;
              imag_value=32707;
            end
    2602  : begin
              real_value= -8477;
              imag_value=31645;
            end
    2603  : begin
              real_value= -14728;
              imag_value=29263;
            end
    2604  : begin
              real_value= -20365;
              imag_value=25661;
            end
    2605  : begin
              real_value= -25154;
              imag_value=20988;
            end
    2606  : begin
              real_value= -28892;
              imag_value=15442;
            end
    2607  : begin
              real_value= -31426;
              imag_value=9253;
            end
    2608  : begin
              real_value= -32651;
              imag_value=2676;
            end
    2609  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    2610  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    2611  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    2612  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    2613  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    2614  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    2615  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    2616  : begin
              real_value= -535;
              imag_value=-32757;
            end
    2617  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    2618  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    2619  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    2620  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    2621  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    2622  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    2623  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    2624  : begin
              real_value= 32721;
              imag_value=1606;
            end
    2625  : begin
              real_value= 31713;
              imag_value=8219;
            end
    2626  : begin
              real_value= 29382;
              imag_value=14489;
            end
    2627  : begin
              real_value= 25826;
              imag_value=20154;
            end
    2628  : begin
              real_value= 21194;
              imag_value=24981;
            end
    2629  : begin
              real_value= 15678;
              imag_value=28766;
            end
    2630  : begin
              real_value= 9508;
              imag_value=31351;
            end
    2631  : begin
              real_value= 2942;
              imag_value=32629;
            end
    2632  : begin
              real_value= -3742;
              imag_value=32547;
            end
    2633  : begin
              real_value= -10275;
              imag_value=31107;
            end
    2634  : begin
              real_value= -16380;
              imag_value=28371;
            end
    2635  : begin
              real_value= -21801;
              imag_value=24453;
            end
    2636  : begin
              real_value= -26314;
              imag_value=19515;
            end
    2637  : begin
              real_value= -29729;
              imag_value=13764;
            end
    2638  : begin
              real_value= -31905;
              imag_value=7438;
            end
    2639  : begin
              real_value= -32750;
              imag_value=802;
            end
    2640  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    2641  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    2642  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    2643  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    2644  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    2645  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    2646  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    2647  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    2648  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    2649  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    2650  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    2651  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    2652  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    2653  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    2654  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    2655  : begin
              real_value= 32575;
              imag_value=3476;
            end
    2656  : begin
              real_value= 31191;
              imag_value=10021;
            end
    2657  : begin
              real_value= 28506;
              imag_value=16148;
            end
    2658  : begin
              real_value= 24630;
              imag_value=21600;
            end
    2659  : begin
              real_value= 19729;
              imag_value=26152;
            end
    2660  : begin
              real_value= 14006;
              imag_value=29615;
            end
    2661  : begin
              real_value= 7699;
              imag_value=31843;
            end
    2662  : begin
              real_value= 1070;
              imag_value=32743;
            end
    2663  : begin
              real_value= -5599;
              imag_value=32278;
            end
    2664  : begin
              real_value= -12039;
              imag_value=30468;
            end
    2665  : begin
              real_value= -17977;
              imag_value=27387;
            end
    2666  : begin
              real_value= -23165;
              imag_value=23165;
            end
    2667  : begin
              real_value= -27387;
              imag_value=17977;
            end
    2668  : begin
              real_value= -30468;
              imag_value=12039;
            end
    2669  : begin
              real_value= -32278;
              imag_value=5599;
            end
    2670  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    2671  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    2672  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    2673  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    2674  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    2675  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    2676  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    2677  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    2678  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    2679  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    2680  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    2681  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    2682  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    2683  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    2684  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    2685  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    2686  : begin
              real_value= 32323;
              imag_value=5336;
            end
    2687  : begin
              real_value= 30565;
              imag_value=11790;
            end
    2688  : begin
              real_value= 27534;
              imag_value=17752;
            end
    2689  : begin
              real_value= 23354;
              imag_value=22974;
            end
    2690  : begin
              real_value= 18200;
              imag_value=27240;
            end
    2691  : begin
              real_value= 12288;
              imag_value=30369;
            end
    2692  : begin
              real_value= 5864;
              imag_value=32231;
            end
    2693  : begin
              real_value= -802;
              imag_value=32750;
            end
    2694  : begin
              real_value= -7438;
              imag_value=31905;
            end
    2695  : begin
              real_value= -13764;
              imag_value=29729;
            end
    2696  : begin
              real_value= -19515;
              imag_value=26314;
            end
    2697  : begin
              real_value= -24453;
              imag_value=21801;
            end
    2698  : begin
              real_value= -28371;
              imag_value=16380;
            end
    2699  : begin
              real_value= -31107;
              imag_value=10275;
            end
    2700  : begin
              real_value= -32547;
              imag_value=3742;
            end
    2701  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    2702  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    2703  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    2704  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    2705  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    2706  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    2707  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    2708  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    2709  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    2710  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    2711  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    2712  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    2713  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    2714  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    2715  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    2716  : begin
              real_value= 32757;
              imag_value=535;
            end
    2717  : begin
              real_value= 31965;
              imag_value=7177;
            end
    2718  : begin
              real_value= 29841;
              imag_value=13520;
            end
    2719  : begin
              real_value= 26472;
              imag_value=19299;
            end
    2720  : begin
              real_value= 22001;
              imag_value=24274;
            end
    2721  : begin
              real_value= 16611;
              imag_value=28236;
            end
    2722  : begin
              real_value= 10529;
              imag_value=31023;
            end
    2723  : begin
              real_value= 4009;
              imag_value=32515;
            end
    2724  : begin
              real_value= -2676;
              imag_value=32651;
            end
    2725  : begin
              real_value= -9253;
              imag_value=31426;
            end
    2726  : begin
              real_value= -15442;
              imag_value=28892;
            end
    2727  : begin
              real_value= -20988;
              imag_value=25154;
            end
    2728  : begin
              real_value= -25661;
              imag_value=20365;
            end
    2729  : begin
              real_value= -29263;
              imag_value=14728;
            end
    2730  : begin
              real_value= -31645;
              imag_value=8477;
            end
    2731  : begin
              real_value= -32707;
              imag_value=1874;
            end
    2732  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    2733  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    2734  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    2735  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    2736  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    2737  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    2738  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    2739  : begin
              real_value= 267;
              imag_value=-32759;
            end
    2740  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    2741  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    2742  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    2743  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    2744  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    2745  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    2746  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    2747  : begin
              real_value= 32673;
              imag_value=2408;
            end
    2748  : begin
              real_value= 31501;
              imag_value=8995;
            end
    2749  : begin
              real_value= 29017;
              imag_value=15206;
            end
    2750  : begin
              real_value= 25324;
              imag_value=20783;
            end
    2751  : begin
              real_value= 20575;
              imag_value=25494;
            end
    2752  : begin
              real_value= 14968;
              imag_value=29142;
            end
    2753  : begin
              real_value= 8737;
              imag_value=31575;
            end
    2754  : begin
              real_value= 2142;
              imag_value=32691;
            end
    2755  : begin
              real_value= -4540;
              imag_value=32445;
            end
    2756  : begin
              real_value= -11036;
              imag_value=30846;
            end
    2757  : begin
              real_value= -17072;
              imag_value=27961;
            end
    2758  : begin
              real_value= -22395;
              imag_value=23911;
            end
    2759  : begin
              real_value= -26784;
              imag_value=18863;
            end
    2760  : begin
              real_value= -30057;
              imag_value=13030;
            end
    2761  : begin
              real_value= -32077;
              imag_value=6654;
            end
    2762  : begin
              real_value= -32760;
              imag_value=0;
            end
    2763  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    2764  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    2765  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    2766  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    2767  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    2768  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    2769  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    2770  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    2771  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    2772  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    2773  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    2774  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    2775  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    2776  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    2777  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    2778  : begin
              real_value= 32481;
              imag_value=4275;
            end
    2779  : begin
              real_value= 30935;
              imag_value=10783;
            end
    2780  : begin
              real_value= 28100;
              imag_value=16842;
            end
    2781  : begin
              real_value= 24092;
              imag_value=22199;
            end
    2782  : begin
              real_value= 19081;
              imag_value=26630;
            end
    2783  : begin
              real_value= 13274;
              imag_value=29950;
            end
    2784  : begin
              real_value= 6915;
              imag_value=32022;
            end
    2785  : begin
              real_value= 267;
              imag_value=32759;
            end
    2786  : begin
              real_value= -6390;
              imag_value=32131;
            end
    2787  : begin
              real_value= -12784;
              imag_value=30163;
            end
    2788  : begin
              real_value= -18644;
              imag_value=26938;
            end
    2789  : begin
              real_value= -23726;
              imag_value=22589;
            end
    2790  : begin
              real_value= -27820;
              imag_value=17299;
            end
    2791  : begin
              real_value= -30755;
              imag_value=11289;
            end
    2792  : begin
              real_value= -32407;
              imag_value=4806;
            end
    2793  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    2794  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    2795  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    2796  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    2797  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    2798  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    2799  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    2800  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    2801  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    2802  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    2803  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    2804  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    2805  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    2806  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    2807  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    2808  : begin
              real_value= 32757;
              imag_value=-535;
            end
    2809  : begin
              real_value= 32183;
              imag_value=6127;
            end
    2810  : begin
              real_value= 30267;
              imag_value=12537;
            end
    2811  : begin
              real_value= 27090;
              imag_value=18423;
            end
    2812  : begin
              real_value= 22782;
              imag_value=23541;
            end
    2813  : begin
              real_value= 17525;
              imag_value=27678;
            end
    2814  : begin
              real_value= 11539;
              imag_value=30661;
            end
    2815  : begin
              real_value= 5071;
              imag_value=32365;
            end
    2816  : begin
              real_value= -1606;
              imag_value=32721;
            end
    2817  : begin
              real_value= -8219;
              imag_value=31713;
            end
    2818  : begin
              real_value= -14489;
              imag_value=29382;
            end
    2819  : begin
              real_value= -20154;
              imag_value=25826;
            end
    2820  : begin
              real_value= -24981;
              imag_value=21194;
            end
    2821  : begin
              real_value= -28766;
              imag_value=15678;
            end
    2822  : begin
              real_value= -31351;
              imag_value=9508;
            end
    2823  : begin
              real_value= -32629;
              imag_value=2942;
            end
    2824  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    2825  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    2826  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    2827  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    2828  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    2829  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    2830  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    2831  : begin
              real_value= -802;
              imag_value=-32750;
            end
    2832  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    2833  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    2834  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    2835  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    2836  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    2837  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    2838  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    2839  : begin
              real_value= 32733;
              imag_value=1338;
            end
    2840  : begin
              real_value= 31779;
              imag_value=7959;
            end
    2841  : begin
              real_value= 29499;
              imag_value=14248;
            end
    2842  : begin
              real_value= 25990;
              imag_value=19943;
            end
    2843  : begin
              real_value= 21399;
              imag_value=24806;
            end
    2844  : begin
              real_value= 15914;
              imag_value=28636;
            end
    2845  : begin
              real_value= 9765;
              imag_value=31271;
            end
    2846  : begin
              real_value= 3210;
              imag_value=32603;
            end
    2847  : begin
              real_value= -3476;
              imag_value=32575;
            end
    2848  : begin
              real_value= -10021;
              imag_value=31191;
            end
    2849  : begin
              real_value= -16148;
              imag_value=28506;
            end
    2850  : begin
              real_value= -21600;
              imag_value=24630;
            end
    2851  : begin
              real_value= -26152;
              imag_value=19729;
            end
    2852  : begin
              real_value= -29615;
              imag_value=14006;
            end
    2853  : begin
              real_value= -31843;
              imag_value=7699;
            end
    2854  : begin
              real_value= -32743;
              imag_value=1070;
            end
    2855  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    2856  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    2857  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    2858  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    2859  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    2860  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    2861  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    2862  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    2863  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    2864  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    2865  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    2866  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    2867  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    2868  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    2869  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    2870  : begin
              real_value= 32603;
              imag_value=3210;
            end
    2871  : begin
              real_value= 31271;
              imag_value=9765;
            end
    2872  : begin
              real_value= 28636;
              imag_value=15914;
            end
    2873  : begin
              real_value= 24806;
              imag_value=21399;
            end
    2874  : begin
              real_value= 19943;
              imag_value=25990;
            end
    2875  : begin
              real_value= 14248;
              imag_value=29499;
            end
    2876  : begin
              real_value= 7959;
              imag_value=31779;
            end
    2877  : begin
              real_value= 1338;
              imag_value=32733;
            end
    2878  : begin
              real_value= -5336;
              imag_value=32323;
            end
    2879  : begin
              real_value= -11790;
              imag_value=30565;
            end
    2880  : begin
              real_value= -17752;
              imag_value=27534;
            end
    2881  : begin
              real_value= -22974;
              imag_value=23354;
            end
    2882  : begin
              real_value= -27240;
              imag_value=18200;
            end
    2883  : begin
              real_value= -30369;
              imag_value=12288;
            end
    2884  : begin
              real_value= -32231;
              imag_value=5864;
            end
    2885  : begin
              real_value= -32750;
              imag_value=-802;
            end
    2886  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    2887  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    2888  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    2889  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    2890  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    2891  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    2892  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    2893  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    2894  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    2895  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    2896  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    2897  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    2898  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    2899  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    2900  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    2901  : begin
              real_value= 32365;
              imag_value=5071;
            end
    2902  : begin
              real_value= 30661;
              imag_value=11539;
            end
    2903  : begin
              real_value= 27678;
              imag_value=17525;
            end
    2904  : begin
              real_value= 23541;
              imag_value=22782;
            end
    2905  : begin
              real_value= 18423;
              imag_value=27090;
            end
    2906  : begin
              real_value= 12537;
              imag_value=30267;
            end
    2907  : begin
              real_value= 6127;
              imag_value=32183;
            end
    2908  : begin
              real_value= -535;
              imag_value=32757;
            end
    2909  : begin
              real_value= -7177;
              imag_value=31965;
            end
    2910  : begin
              real_value= -13520;
              imag_value=29841;
            end
    2911  : begin
              real_value= -19299;
              imag_value=26472;
            end
    2912  : begin
              real_value= -24274;
              imag_value=22001;
            end
    2913  : begin
              real_value= -28236;
              imag_value=16611;
            end
    2914  : begin
              real_value= -31023;
              imag_value=10529;
            end
    2915  : begin
              real_value= -32515;
              imag_value=4009;
            end
    2916  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    2917  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    2918  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    2919  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    2920  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    2921  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    2922  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    2923  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    2924  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    2925  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    2926  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    2927  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    2928  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    2929  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    2930  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    2931  : begin
              real_value= 32759;
              imag_value=267;
            end
    2932  : begin
              real_value= 32022;
              imag_value=6915;
            end
    2933  : begin
              real_value= 29950;
              imag_value=13274;
            end
    2934  : begin
              real_value= 26630;
              imag_value=19081;
            end
    2935  : begin
              real_value= 22199;
              imag_value=24092;
            end
    2936  : begin
              real_value= 16842;
              imag_value=28100;
            end
    2937  : begin
              real_value= 10783;
              imag_value=30935;
            end
    2938  : begin
              real_value= 4275;
              imag_value=32481;
            end
    2939  : begin
              real_value= -2408;
              imag_value=32673;
            end
    2940  : begin
              real_value= -8995;
              imag_value=31501;
            end
    2941  : begin
              real_value= -15206;
              imag_value=29017;
            end
    2942  : begin
              real_value= -20783;
              imag_value=25324;
            end
    2943  : begin
              real_value= -25494;
              imag_value=20575;
            end
    2944  : begin
              real_value= -29142;
              imag_value=14968;
            end
    2945  : begin
              real_value= -31575;
              imag_value=8737;
            end
    2946  : begin
              real_value= -32691;
              imag_value=2142;
            end
    2947  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    2948  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    2949  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    2950  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    2951  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    2952  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    2953  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    2954  : begin
              real_value= 0;
              imag_value=-32760;
            end
    2955  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    2956  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    2957  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    2958  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    2959  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    2960  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    2961  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    2962  : begin
              real_value= 32691;
              imag_value=2142;
            end
    2963  : begin
              real_value= 31575;
              imag_value=8737;
            end
    2964  : begin
              real_value= 29142;
              imag_value=14968;
            end
    2965  : begin
              real_value= 25494;
              imag_value=20575;
            end
    2966  : begin
              real_value= 20783;
              imag_value=25324;
            end
    2967  : begin
              real_value= 15206;
              imag_value=29017;
            end
    2968  : begin
              real_value= 8995;
              imag_value=31501;
            end
    2969  : begin
              real_value= 2408;
              imag_value=32673;
            end
    2970  : begin
              real_value= -4275;
              imag_value=32481;
            end
    2971  : begin
              real_value= -10783;
              imag_value=30935;
            end
    2972  : begin
              real_value= -16842;
              imag_value=28100;
            end
    2973  : begin
              real_value= -22199;
              imag_value=24092;
            end
    2974  : begin
              real_value= -26630;
              imag_value=19081;
            end
    2975  : begin
              real_value= -29950;
              imag_value=13274;
            end
    2976  : begin
              real_value= -32022;
              imag_value=6915;
            end
    2977  : begin
              real_value= -32759;
              imag_value=267;
            end
    2978  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    2979  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    2980  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    2981  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    2982  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    2983  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    2984  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    2985  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    2986  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    2987  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    2988  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    2989  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    2990  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    2991  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    2992  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    2993  : begin
              real_value= 32515;
              imag_value=4009;
            end
    2994  : begin
              real_value= 31023;
              imag_value=10529;
            end
    2995  : begin
              real_value= 28236;
              imag_value=16611;
            end
    2996  : begin
              real_value= 24274;
              imag_value=22001;
            end
    2997  : begin
              real_value= 19299;
              imag_value=26472;
            end
    2998  : begin
              real_value= 13520;
              imag_value=29841;
            end
    2999  : begin
              real_value= 7177;
              imag_value=31965;
            end
    3000  : begin
              real_value= 535;
              imag_value=32757;
            end
    3001  : begin
              real_value= -6127;
              imag_value=32183;
            end
    3002  : begin
              real_value= -12537;
              imag_value=30267;
            end
    3003  : begin
              real_value= -18423;
              imag_value=27090;
            end
    3004  : begin
              real_value= -23541;
              imag_value=22782;
            end
    3005  : begin
              real_value= -27678;
              imag_value=17525;
            end
    3006  : begin
              real_value= -30661;
              imag_value=11539;
            end
    3007  : begin
              real_value= -32365;
              imag_value=5071;
            end
    3008  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    3009  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    3010  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    3011  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    3012  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    3013  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    3014  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    3015  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    3016  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    3017  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    3018  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    3019  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    3020  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    3021  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    3022  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    3023  : begin
              real_value= 32750;
              imag_value=-802;
            end
    3024  : begin
              real_value= 32231;
              imag_value=5864;
            end
    3025  : begin
              real_value= 30369;
              imag_value=12288;
            end
    3026  : begin
              real_value= 27240;
              imag_value=18200;
            end
    3027  : begin
              real_value= 22974;
              imag_value=23354;
            end
    3028  : begin
              real_value= 17752;
              imag_value=27534;
            end
    3029  : begin
              real_value= 11790;
              imag_value=30565;
            end
    3030  : begin
              real_value= 5336;
              imag_value=32323;
            end
    3031  : begin
              real_value= -1338;
              imag_value=32733;
            end
    3032  : begin
              real_value= -7959;
              imag_value=31779;
            end
    3033  : begin
              real_value= -14248;
              imag_value=29499;
            end
    3034  : begin
              real_value= -19943;
              imag_value=25990;
            end
    3035  : begin
              real_value= -24806;
              imag_value=21399;
            end
    3036  : begin
              real_value= -28636;
              imag_value=15914;
            end
    3037  : begin
              real_value= -31271;
              imag_value=9765;
            end
    3038  : begin
              real_value= -32603;
              imag_value=3210;
            end
    3039  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    3040  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    3041  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    3042  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    3043  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    3044  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    3045  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    3046  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    3047  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    3048  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    3049  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    3050  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    3051  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    3052  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    3053  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    3054  : begin
              real_value= 32743;
              imag_value=1070;
            end
    3055  : begin
              real_value= 31843;
              imag_value=7699;
            end
    3056  : begin
              real_value= 29615;
              imag_value=14006;
            end
    3057  : begin
              real_value= 26152;
              imag_value=19729;
            end
    3058  : begin
              real_value= 21600;
              imag_value=24630;
            end
    3059  : begin
              real_value= 16148;
              imag_value=28506;
            end
    3060  : begin
              real_value= 10021;
              imag_value=31191;
            end
    3061  : begin
              real_value= 3476;
              imag_value=32575;
            end
    3062  : begin
              real_value= -3210;
              imag_value=32603;
            end
    3063  : begin
              real_value= -9765;
              imag_value=31271;
            end
    3064  : begin
              real_value= -15914;
              imag_value=28636;
            end
    3065  : begin
              real_value= -21399;
              imag_value=24806;
            end
    3066  : begin
              real_value= -25990;
              imag_value=19943;
            end
    3067  : begin
              real_value= -29499;
              imag_value=14248;
            end
    3068  : begin
              real_value= -31779;
              imag_value=7959;
            end
    3069  : begin
              real_value= -32733;
              imag_value=1338;
            end
    3070  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    3071  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    3072  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    3073  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    3074  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    3075  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    3076  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    3077  : begin
              real_value= 802;
              imag_value=-32750;
            end
    3078  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    3079  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    3080  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    3081  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    3082  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    3083  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    3084  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    3085  : begin
              real_value= 32629;
              imag_value=2942;
            end
    3086  : begin
              real_value= 31351;
              imag_value=9508;
            end
    3087  : begin
              real_value= 28766;
              imag_value=15678;
            end
    3088  : begin
              real_value= 24981;
              imag_value=21194;
            end
    3089  : begin
              real_value= 20154;
              imag_value=25826;
            end
    3090  : begin
              real_value= 14489;
              imag_value=29382;
            end
    3091  : begin
              real_value= 8219;
              imag_value=31713;
            end
    3092  : begin
              real_value= 1606;
              imag_value=32721;
            end
    3093  : begin
              real_value= -5071;
              imag_value=32365;
            end
    3094  : begin
              real_value= -11539;
              imag_value=30661;
            end
    3095  : begin
              real_value= -17525;
              imag_value=27678;
            end
    3096  : begin
              real_value= -22782;
              imag_value=23541;
            end
    3097  : begin
              real_value= -27090;
              imag_value=18423;
            end
    3098  : begin
              real_value= -30267;
              imag_value=12537;
            end
    3099  : begin
              real_value= -32183;
              imag_value=6127;
            end
    3100  : begin
              real_value= -32757;
              imag_value=-535;
            end
    3101  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    3102  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    3103  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    3104  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    3105  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    3106  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    3107  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    3108  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    3109  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    3110  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    3111  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    3112  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    3113  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    3114  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    3115  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    3116  : begin
              real_value= 32407;
              imag_value=4806;
            end
    3117  : begin
              real_value= 30755;
              imag_value=11289;
            end
    3118  : begin
              real_value= 27820;
              imag_value=17299;
            end
    3119  : begin
              real_value= 23726;
              imag_value=22589;
            end
    3120  : begin
              real_value= 18644;
              imag_value=26938;
            end
    3121  : begin
              real_value= 12784;
              imag_value=30163;
            end
    3122  : begin
              real_value= 6390;
              imag_value=32131;
            end
    3123  : begin
              real_value= -267;
              imag_value=32759;
            end
    3124  : begin
              real_value= -6915;
              imag_value=32022;
            end
    3125  : begin
              real_value= -13274;
              imag_value=29950;
            end
    3126  : begin
              real_value= -19081;
              imag_value=26630;
            end
    3127  : begin
              real_value= -24092;
              imag_value=22199;
            end
    3128  : begin
              real_value= -28100;
              imag_value=16842;
            end
    3129  : begin
              real_value= -30935;
              imag_value=10783;
            end
    3130  : begin
              real_value= -32481;
              imag_value=4275;
            end
    3131  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    3132  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    3133  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    3134  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    3135  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    3136  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    3137  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    3138  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    3139  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    3140  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    3141  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    3142  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    3143  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    3144  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    3145  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    3146  : begin
              real_value= 32760;
              imag_value=0;
            end
    3147  : begin
              real_value= 32077;
              imag_value=6654;
            end
    3148  : begin
              real_value= 30057;
              imag_value=13030;
            end
    3149  : begin
              real_value= 26784;
              imag_value=18863;
            end
    3150  : begin
              real_value= 22395;
              imag_value=23911;
            end
    3151  : begin
              real_value= 17072;
              imag_value=27961;
            end
    3152  : begin
              real_value= 11036;
              imag_value=30846;
            end
    3153  : begin
              real_value= 4540;
              imag_value=32445;
            end
    3154  : begin
              real_value= -2142;
              imag_value=32691;
            end
    3155  : begin
              real_value= -8737;
              imag_value=31575;
            end
    3156  : begin
              real_value= -14968;
              imag_value=29142;
            end
    3157  : begin
              real_value= -20575;
              imag_value=25494;
            end
    3158  : begin
              real_value= -25324;
              imag_value=20783;
            end
    3159  : begin
              real_value= -29017;
              imag_value=15206;
            end
    3160  : begin
              real_value= -31501;
              imag_value=8995;
            end
    3161  : begin
              real_value= -32673;
              imag_value=2408;
            end
    3162  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    3163  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    3164  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    3165  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    3166  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    3167  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    3168  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    3169  : begin
              real_value= -267;
              imag_value=-32759;
            end
    3170  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    3171  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    3172  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    3173  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    3174  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    3175  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    3176  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    3177  : begin
              real_value= 32707;
              imag_value=1874;
            end
    3178  : begin
              real_value= 31645;
              imag_value=8477;
            end
    3179  : begin
              real_value= 29263;
              imag_value=14728;
            end
    3180  : begin
              real_value= 25661;
              imag_value=20365;
            end
    3181  : begin
              real_value= 20988;
              imag_value=25154;
            end
    3182  : begin
              real_value= 15442;
              imag_value=28892;
            end
    3183  : begin
              real_value= 9253;
              imag_value=31426;
            end
    3184  : begin
              real_value= 2676;
              imag_value=32651;
            end
    3185  : begin
              real_value= -4009;
              imag_value=32515;
            end
    3186  : begin
              real_value= -10529;
              imag_value=31023;
            end
    3187  : begin
              real_value= -16611;
              imag_value=28236;
            end
    3188  : begin
              real_value= -22001;
              imag_value=24274;
            end
    3189  : begin
              real_value= -26472;
              imag_value=19299;
            end
    3190  : begin
              real_value= -29841;
              imag_value=13520;
            end
    3191  : begin
              real_value= -31965;
              imag_value=7177;
            end
    3192  : begin
              real_value= -32757;
              imag_value=535;
            end
    3193  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    3194  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    3195  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    3196  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    3197  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    3198  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    3199  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    3200  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    3201  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    3202  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    3203  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    3204  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    3205  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    3206  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    3207  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    3208  : begin
              real_value= 32547;
              imag_value=3742;
            end
    3209  : begin
              real_value= 31107;
              imag_value=10275;
            end
    3210  : begin
              real_value= 28371;
              imag_value=16380;
            end
    3211  : begin
              real_value= 24453;
              imag_value=21801;
            end
    3212  : begin
              real_value= 19515;
              imag_value=26314;
            end
    3213  : begin
              real_value= 13764;
              imag_value=29729;
            end
    3214  : begin
              real_value= 7438;
              imag_value=31905;
            end
    3215  : begin
              real_value= 802;
              imag_value=32750;
            end
    3216  : begin
              real_value= -5864;
              imag_value=32231;
            end
    3217  : begin
              real_value= -12288;
              imag_value=30369;
            end
    3218  : begin
              real_value= -18200;
              imag_value=27240;
            end
    3219  : begin
              real_value= -23354;
              imag_value=22974;
            end
    3220  : begin
              real_value= -27534;
              imag_value=17752;
            end
    3221  : begin
              real_value= -30565;
              imag_value=11790;
            end
    3222  : begin
              real_value= -32323;
              imag_value=5336;
            end
    3223  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    3224  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    3225  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    3226  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    3227  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    3228  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    3229  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    3230  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    3231  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    3232  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    3233  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    3234  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    3235  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    3236  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    3237  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    3238  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    3239  : begin
              real_value= 32278;
              imag_value=5599;
            end
    3240  : begin
              real_value= 30468;
              imag_value=12039;
            end
    3241  : begin
              real_value= 27387;
              imag_value=17977;
            end
    3242  : begin
              real_value= 23165;
              imag_value=23165;
            end
    3243  : begin
              real_value= 17977;
              imag_value=27387;
            end
    3244  : begin
              real_value= 12039;
              imag_value=30468;
            end
    3245  : begin
              real_value= 5599;
              imag_value=32278;
            end
    3246  : begin
              real_value= -1070;
              imag_value=32743;
            end
    3247  : begin
              real_value= -7699;
              imag_value=31843;
            end
    3248  : begin
              real_value= -14006;
              imag_value=29615;
            end
    3249  : begin
              real_value= -19729;
              imag_value=26152;
            end
    3250  : begin
              real_value= -24630;
              imag_value=21600;
            end
    3251  : begin
              real_value= -28506;
              imag_value=16148;
            end
    3252  : begin
              real_value= -31191;
              imag_value=10021;
            end
    3253  : begin
              real_value= -32575;
              imag_value=3476;
            end
    3254  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    3255  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    3256  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    3257  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    3258  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    3259  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    3260  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    3261  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    3262  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    3263  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    3264  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    3265  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    3266  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    3267  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    3268  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    3269  : begin
              real_value= 32750;
              imag_value=802;
            end
    3270  : begin
              real_value= 31905;
              imag_value=7438;
            end
    3271  : begin
              real_value= 29729;
              imag_value=13764;
            end
    3272  : begin
              real_value= 26314;
              imag_value=19515;
            end
    3273  : begin
              real_value= 21801;
              imag_value=24453;
            end
    3274  : begin
              real_value= 16380;
              imag_value=28371;
            end
    3275  : begin
              real_value= 10275;
              imag_value=31107;
            end
    3276  : begin
              real_value= 3742;
              imag_value=32547;
            end
    3277  : begin
              real_value= -2942;
              imag_value=32629;
            end
    3278  : begin
              real_value= -9508;
              imag_value=31351;
            end
    3279  : begin
              real_value= -15678;
              imag_value=28766;
            end
    3280  : begin
              real_value= -21194;
              imag_value=24981;
            end
    3281  : begin
              real_value= -25826;
              imag_value=20154;
            end
    3282  : begin
              real_value= -29382;
              imag_value=14489;
            end
    3283  : begin
              real_value= -31713;
              imag_value=8219;
            end
    3284  : begin
              real_value= -32721;
              imag_value=1606;
            end
    3285  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    3286  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    3287  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    3288  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    3289  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    3290  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    3291  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    3292  : begin
              real_value= 535;
              imag_value=-32757;
            end
    3293  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    3294  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    3295  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    3296  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    3297  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    3298  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    3299  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    3300  : begin
              real_value= 32651;
              imag_value=2676;
            end
    3301  : begin
              real_value= 31426;
              imag_value=9253;
            end
    3302  : begin
              real_value= 28892;
              imag_value=15442;
            end
    3303  : begin
              real_value= 25154;
              imag_value=20988;
            end
    3304  : begin
              real_value= 20365;
              imag_value=25661;
            end
    3305  : begin
              real_value= 14728;
              imag_value=29263;
            end
    3306  : begin
              real_value= 8477;
              imag_value=31645;
            end
    3307  : begin
              real_value= 1874;
              imag_value=32707;
            end
    3308  : begin
              real_value= -4806;
              imag_value=32407;
            end
    3309  : begin
              real_value= -11289;
              imag_value=30755;
            end
    3310  : begin
              real_value= -17299;
              imag_value=27820;
            end
    3311  : begin
              real_value= -22589;
              imag_value=23726;
            end
    3312  : begin
              real_value= -26938;
              imag_value=18644;
            end
    3313  : begin
              real_value= -30163;
              imag_value=12784;
            end
    3314  : begin
              real_value= -32131;
              imag_value=6390;
            end
    3315  : begin
              real_value= -32759;
              imag_value=-267;
            end
    3316  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    3317  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    3318  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    3319  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    3320  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    3321  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    3322  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    3323  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    3324  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    3325  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    3326  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    3327  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    3328  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    3329  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    3330  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    3331  : begin
              real_value= 32445;
              imag_value=4540;
            end
    3332  : begin
              real_value= 30846;
              imag_value=11036;
            end
    3333  : begin
              real_value= 27961;
              imag_value=17072;
            end
    3334  : begin
              real_value= 23911;
              imag_value=22395;
            end
    3335  : begin
              real_value= 18863;
              imag_value=26784;
            end
    3336  : begin
              real_value= 13030;
              imag_value=30057;
            end
    3337  : begin
              real_value= 6654;
              imag_value=32077;
            end
    3338  : begin
              real_value= 0;
              imag_value=32760;
            end
    3339  : begin
              real_value= -6654;
              imag_value=32077;
            end
    3340  : begin
              real_value= -13030;
              imag_value=30057;
            end
    3341  : begin
              real_value= -18863;
              imag_value=26784;
            end
    3342  : begin
              real_value= -23911;
              imag_value=22395;
            end
    3343  : begin
              real_value= -27961;
              imag_value=17072;
            end
    3344  : begin
              real_value= -30846;
              imag_value=11036;
            end
    3345  : begin
              real_value= -32445;
              imag_value=4540;
            end
    3346  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    3347  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    3348  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    3349  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    3350  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    3351  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    3352  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    3353  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    3354  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    3355  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    3356  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    3357  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    3358  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    3359  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    3360  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    3361  : begin
              real_value= 32759;
              imag_value=-267;
            end
    3362  : begin
              real_value= 32131;
              imag_value=6390;
            end
    3363  : begin
              real_value= 30163;
              imag_value=12784;
            end
    3364  : begin
              real_value= 26938;
              imag_value=18644;
            end
    3365  : begin
              real_value= 22589;
              imag_value=23726;
            end
    3366  : begin
              real_value= 17299;
              imag_value=27820;
            end
    3367  : begin
              real_value= 11289;
              imag_value=30755;
            end
    3368  : begin
              real_value= 4806;
              imag_value=32407;
            end
    3369  : begin
              real_value= -1874;
              imag_value=32707;
            end
    3370  : begin
              real_value= -8477;
              imag_value=31645;
            end
    3371  : begin
              real_value= -14728;
              imag_value=29263;
            end
    3372  : begin
              real_value= -20365;
              imag_value=25661;
            end
    3373  : begin
              real_value= -25154;
              imag_value=20988;
            end
    3374  : begin
              real_value= -28892;
              imag_value=15442;
            end
    3375  : begin
              real_value= -31426;
              imag_value=9253;
            end
    3376  : begin
              real_value= -32651;
              imag_value=2676;
            end
    3377  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    3378  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    3379  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    3380  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    3381  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    3382  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    3383  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    3384  : begin
              real_value= -535;
              imag_value=-32757;
            end
    3385  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    3386  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    3387  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    3388  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    3389  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    3390  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    3391  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    3392  : begin
              real_value= 32721;
              imag_value=1606;
            end
    3393  : begin
              real_value= 31713;
              imag_value=8219;
            end
    3394  : begin
              real_value= 29382;
              imag_value=14489;
            end
    3395  : begin
              real_value= 25826;
              imag_value=20154;
            end
    3396  : begin
              real_value= 21194;
              imag_value=24981;
            end
    3397  : begin
              real_value= 15678;
              imag_value=28766;
            end
    3398  : begin
              real_value= 9508;
              imag_value=31351;
            end
    3399  : begin
              real_value= 2942;
              imag_value=32629;
            end
    3400  : begin
              real_value= -3742;
              imag_value=32547;
            end
    3401  : begin
              real_value= -10275;
              imag_value=31107;
            end
    3402  : begin
              real_value= -16380;
              imag_value=28371;
            end
    3403  : begin
              real_value= -21801;
              imag_value=24453;
            end
    3404  : begin
              real_value= -26314;
              imag_value=19515;
            end
    3405  : begin
              real_value= -29729;
              imag_value=13764;
            end
    3406  : begin
              real_value= -31905;
              imag_value=7438;
            end
    3407  : begin
              real_value= -32750;
              imag_value=802;
            end
    3408  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    3409  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    3410  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    3411  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    3412  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    3413  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    3414  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    3415  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    3416  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    3417  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    3418  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    3419  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    3420  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    3421  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    3422  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    3423  : begin
              real_value= 32575;
              imag_value=3476;
            end
    3424  : begin
              real_value= 31191;
              imag_value=10021;
            end
    3425  : begin
              real_value= 28506;
              imag_value=16148;
            end
    3426  : begin
              real_value= 24630;
              imag_value=21600;
            end
    3427  : begin
              real_value= 19729;
              imag_value=26152;
            end
    3428  : begin
              real_value= 14006;
              imag_value=29615;
            end
    3429  : begin
              real_value= 7699;
              imag_value=31843;
            end
    3430  : begin
              real_value= 1070;
              imag_value=32743;
            end
    3431  : begin
              real_value= -5599;
              imag_value=32278;
            end
    3432  : begin
              real_value= -12039;
              imag_value=30468;
            end
    3433  : begin
              real_value= -17977;
              imag_value=27387;
            end
    3434  : begin
              real_value= -23165;
              imag_value=23165;
            end
    3435  : begin
              real_value= -27387;
              imag_value=17977;
            end
    3436  : begin
              real_value= -30468;
              imag_value=12039;
            end
    3437  : begin
              real_value= -32278;
              imag_value=5599;
            end
    3438  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    3439  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    3440  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    3441  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    3442  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    3443  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    3444  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    3445  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    3446  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    3447  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    3448  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    3449  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    3450  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    3451  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    3452  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    3453  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    3454  : begin
              real_value= 32323;
              imag_value=5336;
            end
    3455  : begin
              real_value= 30565;
              imag_value=11790;
            end
    3456  : begin
              real_value= 27534;
              imag_value=17752;
            end
    3457  : begin
              real_value= 23354;
              imag_value=22974;
            end
    3458  : begin
              real_value= 18200;
              imag_value=27240;
            end
    3459  : begin
              real_value= 12288;
              imag_value=30369;
            end
    3460  : begin
              real_value= 5864;
              imag_value=32231;
            end
    3461  : begin
              real_value= -802;
              imag_value=32750;
            end
    3462  : begin
              real_value= -7438;
              imag_value=31905;
            end
    3463  : begin
              real_value= -13764;
              imag_value=29729;
            end
    3464  : begin
              real_value= -19515;
              imag_value=26314;
            end
    3465  : begin
              real_value= -24453;
              imag_value=21801;
            end
    3466  : begin
              real_value= -28371;
              imag_value=16380;
            end
    3467  : begin
              real_value= -31107;
              imag_value=10275;
            end
    3468  : begin
              real_value= -32547;
              imag_value=3742;
            end
    3469  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    3470  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    3471  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    3472  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    3473  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    3474  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    3475  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    3476  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    3477  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    3478  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    3479  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    3480  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    3481  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    3482  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    3483  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    3484  : begin
              real_value= 32757;
              imag_value=535;
            end
    3485  : begin
              real_value= 31965;
              imag_value=7177;
            end
    3486  : begin
              real_value= 29841;
              imag_value=13520;
            end
    3487  : begin
              real_value= 26472;
              imag_value=19299;
            end
    3488  : begin
              real_value= 22001;
              imag_value=24274;
            end
    3489  : begin
              real_value= 16611;
              imag_value=28236;
            end
    3490  : begin
              real_value= 10529;
              imag_value=31023;
            end
    3491  : begin
              real_value= 4009;
              imag_value=32515;
            end
    3492  : begin
              real_value= -2676;
              imag_value=32651;
            end
    3493  : begin
              real_value= -9253;
              imag_value=31426;
            end
    3494  : begin
              real_value= -15442;
              imag_value=28892;
            end
    3495  : begin
              real_value= -20988;
              imag_value=25154;
            end
    3496  : begin
              real_value= -25661;
              imag_value=20365;
            end
    3497  : begin
              real_value= -29263;
              imag_value=14728;
            end
    3498  : begin
              real_value= -31645;
              imag_value=8477;
            end
    3499  : begin
              real_value= -32707;
              imag_value=1874;
            end
    3500  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    3501  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    3502  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    3503  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    3504  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    3505  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    3506  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    3507  : begin
              real_value= 267;
              imag_value=-32759;
            end
    3508  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    3509  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    3510  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    3511  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    3512  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    3513  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    3514  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    3515  : begin
              real_value= 32673;
              imag_value=2408;
            end
    3516  : begin
              real_value= 31501;
              imag_value=8995;
            end
    3517  : begin
              real_value= 29017;
              imag_value=15206;
            end
    3518  : begin
              real_value= 25324;
              imag_value=20783;
            end
    3519  : begin
              real_value= 20575;
              imag_value=25494;
            end
    3520  : begin
              real_value= 14968;
              imag_value=29142;
            end
    3521  : begin
              real_value= 8737;
              imag_value=31575;
            end
    3522  : begin
              real_value= 2142;
              imag_value=32691;
            end
    3523  : begin
              real_value= -4540;
              imag_value=32445;
            end
    3524  : begin
              real_value= -11036;
              imag_value=30846;
            end
    3525  : begin
              real_value= -17072;
              imag_value=27961;
            end
    3526  : begin
              real_value= -22395;
              imag_value=23911;
            end
    3527  : begin
              real_value= -26784;
              imag_value=18863;
            end
    3528  : begin
              real_value= -30057;
              imag_value=13030;
            end
    3529  : begin
              real_value= -32077;
              imag_value=6654;
            end
    3530  : begin
              real_value= -32760;
              imag_value=0;
            end
    3531  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    3532  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    3533  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    3534  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    3535  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    3536  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    3537  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    3538  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    3539  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    3540  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    3541  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    3542  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    3543  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    3544  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    3545  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    3546  : begin
              real_value= 32481;
              imag_value=4275;
            end
    3547  : begin
              real_value= 30935;
              imag_value=10783;
            end
    3548  : begin
              real_value= 28100;
              imag_value=16842;
            end
    3549  : begin
              real_value= 24092;
              imag_value=22199;
            end
    3550  : begin
              real_value= 19081;
              imag_value=26630;
            end
    3551  : begin
              real_value= 13274;
              imag_value=29950;
            end
    3552  : begin
              real_value= 6915;
              imag_value=32022;
            end
    3553  : begin
              real_value= 267;
              imag_value=32759;
            end
    3554  : begin
              real_value= -6390;
              imag_value=32131;
            end
    3555  : begin
              real_value= -12784;
              imag_value=30163;
            end
    3556  : begin
              real_value= -18644;
              imag_value=26938;
            end
    3557  : begin
              real_value= -23726;
              imag_value=22589;
            end
    3558  : begin
              real_value= -27820;
              imag_value=17299;
            end
    3559  : begin
              real_value= -30755;
              imag_value=11289;
            end
    3560  : begin
              real_value= -32407;
              imag_value=4806;
            end
    3561  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    3562  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    3563  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    3564  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    3565  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    3566  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    3567  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    3568  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    3569  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    3570  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    3571  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    3572  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    3573  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    3574  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    3575  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    3576  : begin
              real_value= 32757;
              imag_value=-535;
            end
    3577  : begin
              real_value= 32183;
              imag_value=6127;
            end
    3578  : begin
              real_value= 30267;
              imag_value=12537;
            end
    3579  : begin
              real_value= 27090;
              imag_value=18423;
            end
    3580  : begin
              real_value= 22782;
              imag_value=23541;
            end
    3581  : begin
              real_value= 17525;
              imag_value=27678;
            end
    3582  : begin
              real_value= 11539;
              imag_value=30661;
            end
    3583  : begin
              real_value= 5071;
              imag_value=32365;
            end
    3584  : begin
              real_value= -1606;
              imag_value=32721;
            end
    3585  : begin
              real_value= -8219;
              imag_value=31713;
            end
    3586  : begin
              real_value= -14489;
              imag_value=29382;
            end
    3587  : begin
              real_value= -20154;
              imag_value=25826;
            end
    3588  : begin
              real_value= -24981;
              imag_value=21194;
            end
    3589  : begin
              real_value= -28766;
              imag_value=15678;
            end
    3590  : begin
              real_value= -31351;
              imag_value=9508;
            end
    3591  : begin
              real_value= -32629;
              imag_value=2942;
            end
    3592  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    3593  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    3594  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    3595  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    3596  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    3597  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    3598  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    3599  : begin
              real_value= -802;
              imag_value=-32750;
            end
    3600  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    3601  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    3602  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    3603  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    3604  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    3605  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    3606  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    3607  : begin
              real_value= 32733;
              imag_value=1338;
            end
    3608  : begin
              real_value= 31779;
              imag_value=7959;
            end
    3609  : begin
              real_value= 29499;
              imag_value=14248;
            end
    3610  : begin
              real_value= 25990;
              imag_value=19943;
            end
    3611  : begin
              real_value= 21399;
              imag_value=24806;
            end
    3612  : begin
              real_value= 15914;
              imag_value=28636;
            end
    3613  : begin
              real_value= 9765;
              imag_value=31271;
            end
    3614  : begin
              real_value= 3210;
              imag_value=32603;
            end
    3615  : begin
              real_value= -3476;
              imag_value=32575;
            end
    3616  : begin
              real_value= -10021;
              imag_value=31191;
            end
    3617  : begin
              real_value= -16148;
              imag_value=28506;
            end
    3618  : begin
              real_value= -21600;
              imag_value=24630;
            end
    3619  : begin
              real_value= -26152;
              imag_value=19729;
            end
    3620  : begin
              real_value= -29615;
              imag_value=14006;
            end
    3621  : begin
              real_value= -31843;
              imag_value=7699;
            end
    3622  : begin
              real_value= -32743;
              imag_value=1070;
            end
    3623  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    3624  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    3625  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    3626  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    3627  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    3628  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    3629  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    3630  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    3631  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    3632  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    3633  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    3634  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    3635  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    3636  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    3637  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    3638  : begin
              real_value= 32603;
              imag_value=3210;
            end
    3639  : begin
              real_value= 31271;
              imag_value=9765;
            end
    3640  : begin
              real_value= 28636;
              imag_value=15914;
            end
    3641  : begin
              real_value= 24806;
              imag_value=21399;
            end
    3642  : begin
              real_value= 19943;
              imag_value=25990;
            end
    3643  : begin
              real_value= 14248;
              imag_value=29499;
            end
    3644  : begin
              real_value= 7959;
              imag_value=31779;
            end
    3645  : begin
              real_value= 1338;
              imag_value=32733;
            end
    3646  : begin
              real_value= -5336;
              imag_value=32323;
            end
    3647  : begin
              real_value= -11790;
              imag_value=30565;
            end
    3648  : begin
              real_value= -17752;
              imag_value=27534;
            end
    3649  : begin
              real_value= -22974;
              imag_value=23354;
            end
    3650  : begin
              real_value= -27240;
              imag_value=18200;
            end
    3651  : begin
              real_value= -30369;
              imag_value=12288;
            end
    3652  : begin
              real_value= -32231;
              imag_value=5864;
            end
    3653  : begin
              real_value= -32750;
              imag_value=-802;
            end
    3654  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    3655  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    3656  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    3657  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    3658  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    3659  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    3660  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    3661  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    3662  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    3663  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    3664  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    3665  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    3666  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    3667  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    3668  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    3669  : begin
              real_value= 32365;
              imag_value=5071;
            end
    3670  : begin
              real_value= 30661;
              imag_value=11539;
            end
    3671  : begin
              real_value= 27678;
              imag_value=17525;
            end
    3672  : begin
              real_value= 23541;
              imag_value=22782;
            end
    3673  : begin
              real_value= 18423;
              imag_value=27090;
            end
    3674  : begin
              real_value= 12537;
              imag_value=30267;
            end
    3675  : begin
              real_value= 6127;
              imag_value=32183;
            end
    3676  : begin
              real_value= -535;
              imag_value=32757;
            end
    3677  : begin
              real_value= -7177;
              imag_value=31965;
            end
    3678  : begin
              real_value= -13520;
              imag_value=29841;
            end
    3679  : begin
              real_value= -19299;
              imag_value=26472;
            end
    3680  : begin
              real_value= -24274;
              imag_value=22001;
            end
    3681  : begin
              real_value= -28236;
              imag_value=16611;
            end
    3682  : begin
              real_value= -31023;
              imag_value=10529;
            end
    3683  : begin
              real_value= -32515;
              imag_value=4009;
            end
    3684  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    3685  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    3686  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    3687  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    3688  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    3689  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    3690  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    3691  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    3692  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    3693  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    3694  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    3695  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    3696  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    3697  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    3698  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    3699  : begin
              real_value= 32759;
              imag_value=267;
            end
    3700  : begin
              real_value= 32022;
              imag_value=6915;
            end
    3701  : begin
              real_value= 29950;
              imag_value=13274;
            end
    3702  : begin
              real_value= 26630;
              imag_value=19081;
            end
    3703  : begin
              real_value= 22199;
              imag_value=24092;
            end
    3704  : begin
              real_value= 16842;
              imag_value=28100;
            end
    3705  : begin
              real_value= 10783;
              imag_value=30935;
            end
    3706  : begin
              real_value= 4275;
              imag_value=32481;
            end
    3707  : begin
              real_value= -2408;
              imag_value=32673;
            end
    3708  : begin
              real_value= -8995;
              imag_value=31501;
            end
    3709  : begin
              real_value= -15206;
              imag_value=29017;
            end
    3710  : begin
              real_value= -20783;
              imag_value=25324;
            end
    3711  : begin
              real_value= -25494;
              imag_value=20575;
            end
    3712  : begin
              real_value= -29142;
              imag_value=14968;
            end
    3713  : begin
              real_value= -31575;
              imag_value=8737;
            end
    3714  : begin
              real_value= -32691;
              imag_value=2142;
            end
    3715  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    3716  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    3717  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    3718  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    3719  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    3720  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    3721  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    3722  : begin
              real_value= 0;
              imag_value=-32760;
            end
    3723  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    3724  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    3725  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    3726  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    3727  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    3728  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    3729  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    3730  : begin
              real_value= 32691;
              imag_value=2142;
            end
    3731  : begin
              real_value= 31575;
              imag_value=8737;
            end
    3732  : begin
              real_value= 29142;
              imag_value=14968;
            end
    3733  : begin
              real_value= 25494;
              imag_value=20575;
            end
    3734  : begin
              real_value= 20783;
              imag_value=25324;
            end
    3735  : begin
              real_value= 15206;
              imag_value=29017;
            end
    3736  : begin
              real_value= 8995;
              imag_value=31501;
            end
    3737  : begin
              real_value= 2408;
              imag_value=32673;
            end
    3738  : begin
              real_value= -4275;
              imag_value=32481;
            end
    3739  : begin
              real_value= -10783;
              imag_value=30935;
            end
    3740  : begin
              real_value= -16842;
              imag_value=28100;
            end
    3741  : begin
              real_value= -22199;
              imag_value=24092;
            end
    3742  : begin
              real_value= -26630;
              imag_value=19081;
            end
    3743  : begin
              real_value= -29950;
              imag_value=13274;
            end
    3744  : begin
              real_value= -32022;
              imag_value=6915;
            end
    3745  : begin
              real_value= -32759;
              imag_value=267;
            end
    3746  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    3747  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    3748  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    3749  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    3750  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    3751  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    3752  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    3753  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    3754  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    3755  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    3756  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    3757  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    3758  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    3759  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    3760  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    3761  : begin
              real_value= 32515;
              imag_value=4009;
            end
    3762  : begin
              real_value= 31023;
              imag_value=10529;
            end
    3763  : begin
              real_value= 28236;
              imag_value=16611;
            end
    3764  : begin
              real_value= 24274;
              imag_value=22001;
            end
    3765  : begin
              real_value= 19299;
              imag_value=26472;
            end
    3766  : begin
              real_value= 13520;
              imag_value=29841;
            end
    3767  : begin
              real_value= 7177;
              imag_value=31965;
            end
    3768  : begin
              real_value= 535;
              imag_value=32757;
            end
    3769  : begin
              real_value= -6127;
              imag_value=32183;
            end
    3770  : begin
              real_value= -12537;
              imag_value=30267;
            end
    3771  : begin
              real_value= -18423;
              imag_value=27090;
            end
    3772  : begin
              real_value= -23541;
              imag_value=22782;
            end
    3773  : begin
              real_value= -27678;
              imag_value=17525;
            end
    3774  : begin
              real_value= -30661;
              imag_value=11539;
            end
    3775  : begin
              real_value= -32365;
              imag_value=5071;
            end
    3776  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    3777  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    3778  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    3779  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    3780  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    3781  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    3782  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    3783  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    3784  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    3785  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    3786  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    3787  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    3788  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    3789  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    3790  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    3791  : begin
              real_value= 32750;
              imag_value=-802;
            end
    3792  : begin
              real_value= 32231;
              imag_value=5864;
            end
    3793  : begin
              real_value= 30369;
              imag_value=12288;
            end
    3794  : begin
              real_value= 27240;
              imag_value=18200;
            end
    3795  : begin
              real_value= 22974;
              imag_value=23354;
            end
    3796  : begin
              real_value= 17752;
              imag_value=27534;
            end
    3797  : begin
              real_value= 11790;
              imag_value=30565;
            end
    3798  : begin
              real_value= 5336;
              imag_value=32323;
            end
    3799  : begin
              real_value= -1338;
              imag_value=32733;
            end
    3800  : begin
              real_value= -7959;
              imag_value=31779;
            end
    3801  : begin
              real_value= -14248;
              imag_value=29499;
            end
    3802  : begin
              real_value= -19943;
              imag_value=25990;
            end
    3803  : begin
              real_value= -24806;
              imag_value=21399;
            end
    3804  : begin
              real_value= -28636;
              imag_value=15914;
            end
    3805  : begin
              real_value= -31271;
              imag_value=9765;
            end
    3806  : begin
              real_value= -32603;
              imag_value=3210;
            end
    3807  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    3808  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    3809  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    3810  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    3811  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    3812  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    3813  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    3814  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    3815  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    3816  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    3817  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    3818  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    3819  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    3820  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    3821  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    3822  : begin
              real_value= 32743;
              imag_value=1070;
            end
    3823  : begin
              real_value= 31843;
              imag_value=7699;
            end
    3824  : begin
              real_value= 29615;
              imag_value=14006;
            end
    3825  : begin
              real_value= 26152;
              imag_value=19729;
            end
    3826  : begin
              real_value= 21600;
              imag_value=24630;
            end
    3827  : begin
              real_value= 16148;
              imag_value=28506;
            end
    3828  : begin
              real_value= 10021;
              imag_value=31191;
            end
    3829  : begin
              real_value= 3476;
              imag_value=32575;
            end
    3830  : begin
              real_value= -3210;
              imag_value=32603;
            end
    3831  : begin
              real_value= -9765;
              imag_value=31271;
            end
    3832  : begin
              real_value= -15914;
              imag_value=28636;
            end
    3833  : begin
              real_value= -21399;
              imag_value=24806;
            end
    3834  : begin
              real_value= -25990;
              imag_value=19943;
            end
    3835  : begin
              real_value= -29499;
              imag_value=14248;
            end
    3836  : begin
              real_value= -31779;
              imag_value=7959;
            end
    3837  : begin
              real_value= -32733;
              imag_value=1338;
            end
    3838  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    3839  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    3840  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    3841  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    3842  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    3843  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    3844  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    3845  : begin
              real_value= 802;
              imag_value=-32750;
            end
    3846  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    3847  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    3848  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    3849  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    3850  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    3851  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    3852  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    3853  : begin
              real_value= 32629;
              imag_value=2942;
            end
    3854  : begin
              real_value= 31351;
              imag_value=9508;
            end
    3855  : begin
              real_value= 28766;
              imag_value=15678;
            end
    3856  : begin
              real_value= 24981;
              imag_value=21194;
            end
    3857  : begin
              real_value= 20154;
              imag_value=25826;
            end
    3858  : begin
              real_value= 14489;
              imag_value=29382;
            end
    3859  : begin
              real_value= 8219;
              imag_value=31713;
            end
    3860  : begin
              real_value= 1606;
              imag_value=32721;
            end
    3861  : begin
              real_value= -5071;
              imag_value=32365;
            end
    3862  : begin
              real_value= -11539;
              imag_value=30661;
            end
    3863  : begin
              real_value= -17525;
              imag_value=27678;
            end
    3864  : begin
              real_value= -22782;
              imag_value=23541;
            end
    3865  : begin
              real_value= -27090;
              imag_value=18423;
            end
    3866  : begin
              real_value= -30267;
              imag_value=12537;
            end
    3867  : begin
              real_value= -32183;
              imag_value=6127;
            end
    3868  : begin
              real_value= -32757;
              imag_value=-535;
            end
    3869  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    3870  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    3871  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    3872  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    3873  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    3874  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    3875  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    3876  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    3877  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    3878  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    3879  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    3880  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    3881  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    3882  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    3883  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    3884  : begin
              real_value= 32407;
              imag_value=4806;
            end
    3885  : begin
              real_value= 30755;
              imag_value=11289;
            end
    3886  : begin
              real_value= 27820;
              imag_value=17299;
            end
    3887  : begin
              real_value= 23726;
              imag_value=22589;
            end
    3888  : begin
              real_value= 18644;
              imag_value=26938;
            end
    3889  : begin
              real_value= 12784;
              imag_value=30163;
            end
    3890  : begin
              real_value= 6390;
              imag_value=32131;
            end
    3891  : begin
              real_value= -267;
              imag_value=32759;
            end
    3892  : begin
              real_value= -6915;
              imag_value=32022;
            end
    3893  : begin
              real_value= -13274;
              imag_value=29950;
            end
    3894  : begin
              real_value= -19081;
              imag_value=26630;
            end
    3895  : begin
              real_value= -24092;
              imag_value=22199;
            end
    3896  : begin
              real_value= -28100;
              imag_value=16842;
            end
    3897  : begin
              real_value= -30935;
              imag_value=10783;
            end
    3898  : begin
              real_value= -32481;
              imag_value=4275;
            end
    3899  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    3900  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    3901  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    3902  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    3903  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    3904  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    3905  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    3906  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    3907  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    3908  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    3909  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    3910  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    3911  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    3912  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    3913  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    3914  : begin
              real_value= 32760;
              imag_value=0;
            end
    3915  : begin
              real_value= 32077;
              imag_value=6654;
            end
    3916  : begin
              real_value= 30057;
              imag_value=13030;
            end
    3917  : begin
              real_value= 26784;
              imag_value=18863;
            end
    3918  : begin
              real_value= 22395;
              imag_value=23911;
            end
    3919  : begin
              real_value= 17072;
              imag_value=27961;
            end
    3920  : begin
              real_value= 11036;
              imag_value=30846;
            end
    3921  : begin
              real_value= 4540;
              imag_value=32445;
            end
    3922  : begin
              real_value= -2142;
              imag_value=32691;
            end
    3923  : begin
              real_value= -8737;
              imag_value=31575;
            end
    3924  : begin
              real_value= -14968;
              imag_value=29142;
            end
    3925  : begin
              real_value= -20575;
              imag_value=25494;
            end
    3926  : begin
              real_value= -25324;
              imag_value=20783;
            end
    3927  : begin
              real_value= -29017;
              imag_value=15206;
            end
    3928  : begin
              real_value= -31501;
              imag_value=8995;
            end
    3929  : begin
              real_value= -32673;
              imag_value=2408;
            end
    3930  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    3931  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    3932  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    3933  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    3934  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    3935  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    3936  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    3937  : begin
              real_value= -267;
              imag_value=-32759;
            end
    3938  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    3939  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    3940  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    3941  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    3942  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    3943  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    3944  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    3945  : begin
              real_value= 32707;
              imag_value=1874;
            end
    3946  : begin
              real_value= 31645;
              imag_value=8477;
            end
    3947  : begin
              real_value= 29263;
              imag_value=14728;
            end
    3948  : begin
              real_value= 25661;
              imag_value=20365;
            end
    3949  : begin
              real_value= 20988;
              imag_value=25154;
            end
    3950  : begin
              real_value= 15442;
              imag_value=28892;
            end
    3951  : begin
              real_value= 9253;
              imag_value=31426;
            end
    3952  : begin
              real_value= 2676;
              imag_value=32651;
            end
    3953  : begin
              real_value= -4009;
              imag_value=32515;
            end
    3954  : begin
              real_value= -10529;
              imag_value=31023;
            end
    3955  : begin
              real_value= -16611;
              imag_value=28236;
            end
    3956  : begin
              real_value= -22001;
              imag_value=24274;
            end
    3957  : begin
              real_value= -26472;
              imag_value=19299;
            end
    3958  : begin
              real_value= -29841;
              imag_value=13520;
            end
    3959  : begin
              real_value= -31965;
              imag_value=7177;
            end
    3960  : begin
              real_value= -32757;
              imag_value=535;
            end
    3961  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    3962  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    3963  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    3964  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    3965  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    3966  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    3967  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    3968  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    3969  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    3970  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    3971  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    3972  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    3973  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    3974  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    3975  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    3976  : begin
              real_value= 32547;
              imag_value=3742;
            end
    3977  : begin
              real_value= 31107;
              imag_value=10275;
            end
    3978  : begin
              real_value= 28371;
              imag_value=16380;
            end
    3979  : begin
              real_value= 24453;
              imag_value=21801;
            end
    3980  : begin
              real_value= 19515;
              imag_value=26314;
            end
    3981  : begin
              real_value= 13764;
              imag_value=29729;
            end
    3982  : begin
              real_value= 7438;
              imag_value=31905;
            end
    3983  : begin
              real_value= 802;
              imag_value=32750;
            end
    3984  : begin
              real_value= -5864;
              imag_value=32231;
            end
    3985  : begin
              real_value= -12288;
              imag_value=30369;
            end
    3986  : begin
              real_value= -18200;
              imag_value=27240;
            end
    3987  : begin
              real_value= -23354;
              imag_value=22974;
            end
    3988  : begin
              real_value= -27534;
              imag_value=17752;
            end
    3989  : begin
              real_value= -30565;
              imag_value=11790;
            end
    3990  : begin
              real_value= -32323;
              imag_value=5336;
            end
    3991  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    3992  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    3993  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    3994  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    3995  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    3996  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    3997  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    3998  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    3999  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    4000  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    4001  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    4002  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    4003  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    4004  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    4005  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    4006  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    4007  : begin
              real_value= 32278;
              imag_value=5599;
            end
    4008  : begin
              real_value= 30468;
              imag_value=12039;
            end
    4009  : begin
              real_value= 27387;
              imag_value=17977;
            end
    4010  : begin
              real_value= 23165;
              imag_value=23165;
            end
    4011  : begin
              real_value= 17977;
              imag_value=27387;
            end
    4012  : begin
              real_value= 12039;
              imag_value=30468;
            end
    4013  : begin
              real_value= 5599;
              imag_value=32278;
            end
    4014  : begin
              real_value= -1070;
              imag_value=32743;
            end
    4015  : begin
              real_value= -7699;
              imag_value=31843;
            end
    4016  : begin
              real_value= -14006;
              imag_value=29615;
            end
    4017  : begin
              real_value= -19729;
              imag_value=26152;
            end
    4018  : begin
              real_value= -24630;
              imag_value=21600;
            end
    4019  : begin
              real_value= -28506;
              imag_value=16148;
            end
    4020  : begin
              real_value= -31191;
              imag_value=10021;
            end
    4021  : begin
              real_value= -32575;
              imag_value=3476;
            end
    4022  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    4023  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    4024  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    4025  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    4026  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    4027  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    4028  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    4029  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    4030  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    4031  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    4032  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    4033  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    4034  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    4035  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    4036  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    4037  : begin
              real_value= 32750;
              imag_value=802;
            end
    4038  : begin
              real_value= 31905;
              imag_value=7438;
            end
    4039  : begin
              real_value= 29729;
              imag_value=13764;
            end
    4040  : begin
              real_value= 26314;
              imag_value=19515;
            end
    4041  : begin
              real_value= 21801;
              imag_value=24453;
            end
    4042  : begin
              real_value= 16380;
              imag_value=28371;
            end
    4043  : begin
              real_value= 10275;
              imag_value=31107;
            end
    4044  : begin
              real_value= 3742;
              imag_value=32547;
            end
    4045  : begin
              real_value= -2942;
              imag_value=32629;
            end
    4046  : begin
              real_value= -9508;
              imag_value=31351;
            end
    4047  : begin
              real_value= -15678;
              imag_value=28766;
            end
    4048  : begin
              real_value= -21194;
              imag_value=24981;
            end
    4049  : begin
              real_value= -25826;
              imag_value=20154;
            end
    4050  : begin
              real_value= -29382;
              imag_value=14489;
            end
    4051  : begin
              real_value= -31713;
              imag_value=8219;
            end
    4052  : begin
              real_value= -32721;
              imag_value=1606;
            end
    4053  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    4054  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    4055  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    4056  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    4057  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    4058  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    4059  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    4060  : begin
              real_value= 535;
              imag_value=-32757;
            end
    4061  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    4062  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    4063  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    4064  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    4065  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    4066  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    4067  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    4068  : begin
              real_value= 32651;
              imag_value=2676;
            end
    4069  : begin
              real_value= 31426;
              imag_value=9253;
            end
    4070  : begin
              real_value= 28892;
              imag_value=15442;
            end
    4071  : begin
              real_value= 25154;
              imag_value=20988;
            end
    4072  : begin
              real_value= 20365;
              imag_value=25661;
            end
    4073  : begin
              real_value= 14728;
              imag_value=29263;
            end
    4074  : begin
              real_value= 8477;
              imag_value=31645;
            end
    4075  : begin
              real_value= 1874;
              imag_value=32707;
            end
    4076  : begin
              real_value= -4806;
              imag_value=32407;
            end
    4077  : begin
              real_value= -11289;
              imag_value=30755;
            end
    4078  : begin
              real_value= -17299;
              imag_value=27820;
            end
    4079  : begin
              real_value= -22589;
              imag_value=23726;
            end
    4080  : begin
              real_value= -26938;
              imag_value=18644;
            end
    4081  : begin
              real_value= -30163;
              imag_value=12784;
            end
    4082  : begin
              real_value= -32131;
              imag_value=6390;
            end
    4083  : begin
              real_value= -32759;
              imag_value=-267;
            end
    4084  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    4085  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    4086  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    4087  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    4088  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    4089  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    4090  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    4091  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    4092  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    4093  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    4094  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    4095  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    4096  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    4097  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    4098  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    4099  : begin
              real_value= 32445;
              imag_value=4540;
            end
    4100  : begin
              real_value= 30846;
              imag_value=11036;
            end
    4101  : begin
              real_value= 27961;
              imag_value=17072;
            end
    4102  : begin
              real_value= 23911;
              imag_value=22395;
            end
    4103  : begin
              real_value= 18863;
              imag_value=26784;
            end
    4104  : begin
              real_value= 13030;
              imag_value=30057;
            end
    4105  : begin
              real_value= 6654;
              imag_value=32077;
            end
    4106  : begin
              real_value= 0;
              imag_value=32760;
            end
    4107  : begin
              real_value= -6654;
              imag_value=32077;
            end
    4108  : begin
              real_value= -13030;
              imag_value=30057;
            end
    4109  : begin
              real_value= -18863;
              imag_value=26784;
            end
    4110  : begin
              real_value= -23911;
              imag_value=22395;
            end
    4111  : begin
              real_value= -27961;
              imag_value=17072;
            end
    4112  : begin
              real_value= -30846;
              imag_value=11036;
            end
    4113  : begin
              real_value= -32445;
              imag_value=4540;
            end
    4114  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    4115  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    4116  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    4117  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    4118  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    4119  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    4120  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    4121  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    4122  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    4123  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    4124  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    4125  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    4126  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    4127  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    4128  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    4129  : begin
              real_value= 32759;
              imag_value=-267;
            end
    4130  : begin
              real_value= 32131;
              imag_value=6390;
            end
    4131  : begin
              real_value= 30163;
              imag_value=12784;
            end
    4132  : begin
              real_value= 26938;
              imag_value=18644;
            end
    4133  : begin
              real_value= 22589;
              imag_value=23726;
            end
    4134  : begin
              real_value= 17299;
              imag_value=27820;
            end
    4135  : begin
              real_value= 11289;
              imag_value=30755;
            end
    4136  : begin
              real_value= 4806;
              imag_value=32407;
            end
    4137  : begin
              real_value= -1874;
              imag_value=32707;
            end
    4138  : begin
              real_value= -8477;
              imag_value=31645;
            end
    4139  : begin
              real_value= -14728;
              imag_value=29263;
            end
    4140  : begin
              real_value= -20365;
              imag_value=25661;
            end
    4141  : begin
              real_value= -25154;
              imag_value=20988;
            end
    4142  : begin
              real_value= -28892;
              imag_value=15442;
            end
    4143  : begin
              real_value= -31426;
              imag_value=9253;
            end
    4144  : begin
              real_value= -32651;
              imag_value=2676;
            end
    4145  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    4146  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    4147  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    4148  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    4149  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    4150  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    4151  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    4152  : begin
              real_value= -535;
              imag_value=-32757;
            end
    4153  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    4154  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    4155  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    4156  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    4157  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    4158  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    4159  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    4160  : begin
              real_value= 32721;
              imag_value=1606;
            end
    4161  : begin
              real_value= 31713;
              imag_value=8219;
            end
    4162  : begin
              real_value= 29382;
              imag_value=14489;
            end
    4163  : begin
              real_value= 25826;
              imag_value=20154;
            end
    4164  : begin
              real_value= 21194;
              imag_value=24981;
            end
    4165  : begin
              real_value= 15678;
              imag_value=28766;
            end
    4166  : begin
              real_value= 9508;
              imag_value=31351;
            end
    4167  : begin
              real_value= 2942;
              imag_value=32629;
            end
    4168  : begin
              real_value= -3742;
              imag_value=32547;
            end
    4169  : begin
              real_value= -10275;
              imag_value=31107;
            end
    4170  : begin
              real_value= -16380;
              imag_value=28371;
            end
    4171  : begin
              real_value= -21801;
              imag_value=24453;
            end
    4172  : begin
              real_value= -26314;
              imag_value=19515;
            end
    4173  : begin
              real_value= -29729;
              imag_value=13764;
            end
    4174  : begin
              real_value= -31905;
              imag_value=7438;
            end
    4175  : begin
              real_value= -32750;
              imag_value=802;
            end
    4176  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    4177  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    4178  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    4179  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    4180  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    4181  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    4182  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    4183  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    4184  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    4185  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    4186  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    4187  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    4188  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    4189  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    4190  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    4191  : begin
              real_value= 32575;
              imag_value=3476;
            end
    4192  : begin
              real_value= 31191;
              imag_value=10021;
            end
    4193  : begin
              real_value= 28506;
              imag_value=16148;
            end
    4194  : begin
              real_value= 24630;
              imag_value=21600;
            end
    4195  : begin
              real_value= 19729;
              imag_value=26152;
            end
    4196  : begin
              real_value= 14006;
              imag_value=29615;
            end
    4197  : begin
              real_value= 7699;
              imag_value=31843;
            end
    4198  : begin
              real_value= 1070;
              imag_value=32743;
            end
    4199  : begin
              real_value= -5599;
              imag_value=32278;
            end
    4200  : begin
              real_value= -12039;
              imag_value=30468;
            end
    4201  : begin
              real_value= -17977;
              imag_value=27387;
            end
    4202  : begin
              real_value= -23165;
              imag_value=23165;
            end
    4203  : begin
              real_value= -27387;
              imag_value=17977;
            end
    4204  : begin
              real_value= -30468;
              imag_value=12039;
            end
    4205  : begin
              real_value= -32278;
              imag_value=5599;
            end
    4206  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    4207  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    4208  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    4209  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    4210  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    4211  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    4212  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    4213  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    4214  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    4215  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    4216  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    4217  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    4218  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    4219  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    4220  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    4221  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    4222  : begin
              real_value= 32323;
              imag_value=5336;
            end
    4223  : begin
              real_value= 30565;
              imag_value=11790;
            end
    4224  : begin
              real_value= 27534;
              imag_value=17752;
            end
    4225  : begin
              real_value= 23354;
              imag_value=22974;
            end
    4226  : begin
              real_value= 18200;
              imag_value=27240;
            end
    4227  : begin
              real_value= 12288;
              imag_value=30369;
            end
    4228  : begin
              real_value= 5864;
              imag_value=32231;
            end
    4229  : begin
              real_value= -802;
              imag_value=32750;
            end
    4230  : begin
              real_value= -7438;
              imag_value=31905;
            end
    4231  : begin
              real_value= -13764;
              imag_value=29729;
            end
    4232  : begin
              real_value= -19515;
              imag_value=26314;
            end
    4233  : begin
              real_value= -24453;
              imag_value=21801;
            end
    4234  : begin
              real_value= -28371;
              imag_value=16380;
            end
    4235  : begin
              real_value= -31107;
              imag_value=10275;
            end
    4236  : begin
              real_value= -32547;
              imag_value=3742;
            end
    4237  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    4238  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    4239  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    4240  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    4241  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    4242  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    4243  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    4244  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    4245  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    4246  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    4247  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    4248  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    4249  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    4250  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    4251  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    4252  : begin
              real_value= 32757;
              imag_value=535;
            end
    4253  : begin
              real_value= 31965;
              imag_value=7177;
            end
    4254  : begin
              real_value= 29841;
              imag_value=13520;
            end
    4255  : begin
              real_value= 26472;
              imag_value=19299;
            end
    4256  : begin
              real_value= 22001;
              imag_value=24274;
            end
    4257  : begin
              real_value= 16611;
              imag_value=28236;
            end
    4258  : begin
              real_value= 10529;
              imag_value=31023;
            end
    4259  : begin
              real_value= 4009;
              imag_value=32515;
            end
    4260  : begin
              real_value= -2676;
              imag_value=32651;
            end
    4261  : begin
              real_value= -9253;
              imag_value=31426;
            end
    4262  : begin
              real_value= -15442;
              imag_value=28892;
            end
    4263  : begin
              real_value= -20988;
              imag_value=25154;
            end
    4264  : begin
              real_value= -25661;
              imag_value=20365;
            end
    4265  : begin
              real_value= -29263;
              imag_value=14728;
            end
    4266  : begin
              real_value= -31645;
              imag_value=8477;
            end
    4267  : begin
              real_value= -32707;
              imag_value=1874;
            end
    4268  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    4269  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    4270  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    4271  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    4272  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    4273  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    4274  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    4275  : begin
              real_value= 267;
              imag_value=-32759;
            end
    4276  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    4277  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    4278  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    4279  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    4280  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    4281  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    4282  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    4283  : begin
              real_value= 32673;
              imag_value=2408;
            end
    4284  : begin
              real_value= 31501;
              imag_value=8995;
            end
    4285  : begin
              real_value= 29017;
              imag_value=15206;
            end
    4286  : begin
              real_value= 25324;
              imag_value=20783;
            end
    4287  : begin
              real_value= 20575;
              imag_value=25494;
            end
    4288  : begin
              real_value= 14968;
              imag_value=29142;
            end
    4289  : begin
              real_value= 8737;
              imag_value=31575;
            end
    4290  : begin
              real_value= 2142;
              imag_value=32691;
            end
    4291  : begin
              real_value= -4540;
              imag_value=32445;
            end
    4292  : begin
              real_value= -11036;
              imag_value=30846;
            end
    4293  : begin
              real_value= -17072;
              imag_value=27961;
            end
    4294  : begin
              real_value= -22395;
              imag_value=23911;
            end
    4295  : begin
              real_value= -26784;
              imag_value=18863;
            end
    4296  : begin
              real_value= -30057;
              imag_value=13030;
            end
    4297  : begin
              real_value= -32077;
              imag_value=6654;
            end
    4298  : begin
              real_value= -32760;
              imag_value=0;
            end
    4299  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    4300  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    4301  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    4302  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    4303  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    4304  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    4305  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    4306  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    4307  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    4308  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    4309  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    4310  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    4311  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    4312  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    4313  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    4314  : begin
              real_value= 32481;
              imag_value=4275;
            end
    4315  : begin
              real_value= 30935;
              imag_value=10783;
            end
    4316  : begin
              real_value= 28100;
              imag_value=16842;
            end
    4317  : begin
              real_value= 24092;
              imag_value=22199;
            end
    4318  : begin
              real_value= 19081;
              imag_value=26630;
            end
    4319  : begin
              real_value= 13274;
              imag_value=29950;
            end
    4320  : begin
              real_value= 6915;
              imag_value=32022;
            end
    4321  : begin
              real_value= 267;
              imag_value=32759;
            end
    4322  : begin
              real_value= -6390;
              imag_value=32131;
            end
    4323  : begin
              real_value= -12784;
              imag_value=30163;
            end
    4324  : begin
              real_value= -18644;
              imag_value=26938;
            end
    4325  : begin
              real_value= -23726;
              imag_value=22589;
            end
    4326  : begin
              real_value= -27820;
              imag_value=17299;
            end
    4327  : begin
              real_value= -30755;
              imag_value=11289;
            end
    4328  : begin
              real_value= -32407;
              imag_value=4806;
            end
    4329  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    4330  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    4331  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    4332  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    4333  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    4334  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    4335  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    4336  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    4337  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    4338  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    4339  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    4340  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    4341  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    4342  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    4343  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    4344  : begin
              real_value= 32757;
              imag_value=-535;
            end
    4345  : begin
              real_value= 32183;
              imag_value=6127;
            end
    4346  : begin
              real_value= 30267;
              imag_value=12537;
            end
    4347  : begin
              real_value= 27090;
              imag_value=18423;
            end
    4348  : begin
              real_value= 22782;
              imag_value=23541;
            end
    4349  : begin
              real_value= 17525;
              imag_value=27678;
            end
    4350  : begin
              real_value= 11539;
              imag_value=30661;
            end
    4351  : begin
              real_value= 5071;
              imag_value=32365;
            end
    4352  : begin
              real_value= -1606;
              imag_value=32721;
            end
    4353  : begin
              real_value= -8219;
              imag_value=31713;
            end
    4354  : begin
              real_value= -14489;
              imag_value=29382;
            end
    4355  : begin
              real_value= -20154;
              imag_value=25826;
            end
    4356  : begin
              real_value= -24981;
              imag_value=21194;
            end
    4357  : begin
              real_value= -28766;
              imag_value=15678;
            end
    4358  : begin
              real_value= -31351;
              imag_value=9508;
            end
    4359  : begin
              real_value= -32629;
              imag_value=2942;
            end
    4360  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    4361  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    4362  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    4363  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    4364  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    4365  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    4366  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    4367  : begin
              real_value= -802;
              imag_value=-32750;
            end
    4368  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    4369  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    4370  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    4371  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    4372  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    4373  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    4374  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    4375  : begin
              real_value= 32733;
              imag_value=1338;
            end
    4376  : begin
              real_value= 31779;
              imag_value=7959;
            end
    4377  : begin
              real_value= 29499;
              imag_value=14248;
            end
    4378  : begin
              real_value= 25990;
              imag_value=19943;
            end
    4379  : begin
              real_value= 21399;
              imag_value=24806;
            end
    4380  : begin
              real_value= 15914;
              imag_value=28636;
            end
    4381  : begin
              real_value= 9765;
              imag_value=31271;
            end
    4382  : begin
              real_value= 3210;
              imag_value=32603;
            end
    4383  : begin
              real_value= -3476;
              imag_value=32575;
            end
    4384  : begin
              real_value= -10021;
              imag_value=31191;
            end
    4385  : begin
              real_value= -16148;
              imag_value=28506;
            end
    4386  : begin
              real_value= -21600;
              imag_value=24630;
            end
    4387  : begin
              real_value= -26152;
              imag_value=19729;
            end
    4388  : begin
              real_value= -29615;
              imag_value=14006;
            end
    4389  : begin
              real_value= -31843;
              imag_value=7699;
            end
    4390  : begin
              real_value= -32743;
              imag_value=1070;
            end
    4391  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    4392  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    4393  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    4394  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    4395  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    4396  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    4397  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    4398  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    4399  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    4400  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    4401  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    4402  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    4403  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    4404  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    4405  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    4406  : begin
              real_value= 32603;
              imag_value=3210;
            end
    4407  : begin
              real_value= 31271;
              imag_value=9765;
            end
    4408  : begin
              real_value= 28636;
              imag_value=15914;
            end
    4409  : begin
              real_value= 24806;
              imag_value=21399;
            end
    4410  : begin
              real_value= 19943;
              imag_value=25990;
            end
    4411  : begin
              real_value= 14248;
              imag_value=29499;
            end
    4412  : begin
              real_value= 7959;
              imag_value=31779;
            end
    4413  : begin
              real_value= 1338;
              imag_value=32733;
            end
    4414  : begin
              real_value= -5336;
              imag_value=32323;
            end
    4415  : begin
              real_value= -11790;
              imag_value=30565;
            end
    4416  : begin
              real_value= -17752;
              imag_value=27534;
            end
    4417  : begin
              real_value= -22974;
              imag_value=23354;
            end
    4418  : begin
              real_value= -27240;
              imag_value=18200;
            end
    4419  : begin
              real_value= -30369;
              imag_value=12288;
            end
    4420  : begin
              real_value= -32231;
              imag_value=5864;
            end
    4421  : begin
              real_value= -32750;
              imag_value=-802;
            end
    4422  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    4423  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    4424  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    4425  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    4426  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    4427  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    4428  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    4429  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    4430  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    4431  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    4432  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    4433  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    4434  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    4435  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    4436  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    4437  : begin
              real_value= 32365;
              imag_value=5071;
            end
    4438  : begin
              real_value= 30661;
              imag_value=11539;
            end
    4439  : begin
              real_value= 27678;
              imag_value=17525;
            end
    4440  : begin
              real_value= 23541;
              imag_value=22782;
            end
    4441  : begin
              real_value= 18423;
              imag_value=27090;
            end
    4442  : begin
              real_value= 12537;
              imag_value=30267;
            end
    4443  : begin
              real_value= 6127;
              imag_value=32183;
            end
    4444  : begin
              real_value= -535;
              imag_value=32757;
            end
    4445  : begin
              real_value= -7177;
              imag_value=31965;
            end
    4446  : begin
              real_value= -13520;
              imag_value=29841;
            end
    4447  : begin
              real_value= -19299;
              imag_value=26472;
            end
    4448  : begin
              real_value= -24274;
              imag_value=22001;
            end
    4449  : begin
              real_value= -28236;
              imag_value=16611;
            end
    4450  : begin
              real_value= -31023;
              imag_value=10529;
            end
    4451  : begin
              real_value= -32515;
              imag_value=4009;
            end
    4452  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    4453  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    4454  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    4455  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    4456  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    4457  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    4458  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    4459  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    4460  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    4461  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    4462  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    4463  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    4464  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    4465  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    4466  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    4467  : begin
              real_value= 32759;
              imag_value=267;
            end
    4468  : begin
              real_value= 32022;
              imag_value=6915;
            end
    4469  : begin
              real_value= 29950;
              imag_value=13274;
            end
    4470  : begin
              real_value= 26630;
              imag_value=19081;
            end
    4471  : begin
              real_value= 22199;
              imag_value=24092;
            end
    4472  : begin
              real_value= 16842;
              imag_value=28100;
            end
    4473  : begin
              real_value= 10783;
              imag_value=30935;
            end
    4474  : begin
              real_value= 4275;
              imag_value=32481;
            end
    4475  : begin
              real_value= -2408;
              imag_value=32673;
            end
    4476  : begin
              real_value= -8995;
              imag_value=31501;
            end
    4477  : begin
              real_value= -15206;
              imag_value=29017;
            end
    4478  : begin
              real_value= -20783;
              imag_value=25324;
            end
    4479  : begin
              real_value= -25494;
              imag_value=20575;
            end
    4480  : begin
              real_value= -29142;
              imag_value=14968;
            end
    4481  : begin
              real_value= -31575;
              imag_value=8737;
            end
    4482  : begin
              real_value= -32691;
              imag_value=2142;
            end
    4483  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    4484  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    4485  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    4486  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    4487  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    4488  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    4489  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    4490  : begin
              real_value= 0;
              imag_value=-32760;
            end
    4491  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    4492  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    4493  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    4494  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    4495  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    4496  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    4497  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    4498  : begin
              real_value= 32691;
              imag_value=2142;
            end
    4499  : begin
              real_value= 31575;
              imag_value=8737;
            end
    4500  : begin
              real_value= 29142;
              imag_value=14968;
            end
    4501  : begin
              real_value= 25494;
              imag_value=20575;
            end
    4502  : begin
              real_value= 20783;
              imag_value=25324;
            end
    4503  : begin
              real_value= 15206;
              imag_value=29017;
            end
    4504  : begin
              real_value= 8995;
              imag_value=31501;
            end
    4505  : begin
              real_value= 2408;
              imag_value=32673;
            end
    4506  : begin
              real_value= -4275;
              imag_value=32481;
            end
    4507  : begin
              real_value= -10783;
              imag_value=30935;
            end
    4508  : begin
              real_value= -16842;
              imag_value=28100;
            end
    4509  : begin
              real_value= -22199;
              imag_value=24092;
            end
    4510  : begin
              real_value= -26630;
              imag_value=19081;
            end
    4511  : begin
              real_value= -29950;
              imag_value=13274;
            end
    4512  : begin
              real_value= -32022;
              imag_value=6915;
            end
    4513  : begin
              real_value= -32759;
              imag_value=267;
            end
    4514  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    4515  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    4516  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    4517  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    4518  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    4519  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    4520  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    4521  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    4522  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    4523  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    4524  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    4525  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    4526  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    4527  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    4528  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    4529  : begin
              real_value= 32515;
              imag_value=4009;
            end
    4530  : begin
              real_value= 31023;
              imag_value=10529;
            end
    4531  : begin
              real_value= 28236;
              imag_value=16611;
            end
    4532  : begin
              real_value= 24274;
              imag_value=22001;
            end
    4533  : begin
              real_value= 19299;
              imag_value=26472;
            end
    4534  : begin
              real_value= 13520;
              imag_value=29841;
            end
    4535  : begin
              real_value= 7177;
              imag_value=31965;
            end
    4536  : begin
              real_value= 535;
              imag_value=32757;
            end
    4537  : begin
              real_value= -6127;
              imag_value=32183;
            end
    4538  : begin
              real_value= -12537;
              imag_value=30267;
            end
    4539  : begin
              real_value= -18423;
              imag_value=27090;
            end
    4540  : begin
              real_value= -23541;
              imag_value=22782;
            end
    4541  : begin
              real_value= -27678;
              imag_value=17525;
            end
    4542  : begin
              real_value= -30661;
              imag_value=11539;
            end
    4543  : begin
              real_value= -32365;
              imag_value=5071;
            end
    4544  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    4545  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    4546  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    4547  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    4548  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    4549  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    4550  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    4551  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    4552  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    4553  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    4554  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    4555  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    4556  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    4557  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    4558  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    4559  : begin
              real_value= 32750;
              imag_value=-802;
            end
    4560  : begin
              real_value= 32231;
              imag_value=5864;
            end
    4561  : begin
              real_value= 30369;
              imag_value=12288;
            end
    4562  : begin
              real_value= 27240;
              imag_value=18200;
            end
    4563  : begin
              real_value= 22974;
              imag_value=23354;
            end
    4564  : begin
              real_value= 17752;
              imag_value=27534;
            end
    4565  : begin
              real_value= 11790;
              imag_value=30565;
            end
    4566  : begin
              real_value= 5336;
              imag_value=32323;
            end
    4567  : begin
              real_value= -1338;
              imag_value=32733;
            end
    4568  : begin
              real_value= -7959;
              imag_value=31779;
            end
    4569  : begin
              real_value= -14248;
              imag_value=29499;
            end
    4570  : begin
              real_value= -19943;
              imag_value=25990;
            end
    4571  : begin
              real_value= -24806;
              imag_value=21399;
            end
    4572  : begin
              real_value= -28636;
              imag_value=15914;
            end
    4573  : begin
              real_value= -31271;
              imag_value=9765;
            end
    4574  : begin
              real_value= -32603;
              imag_value=3210;
            end
    4575  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    4576  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    4577  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    4578  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    4579  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    4580  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    4581  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    4582  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    4583  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    4584  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    4585  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    4586  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    4587  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    4588  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    4589  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    4590  : begin
              real_value= 32743;
              imag_value=1070;
            end
    4591  : begin
              real_value= 31843;
              imag_value=7699;
            end
    4592  : begin
              real_value= 29615;
              imag_value=14006;
            end
    4593  : begin
              real_value= 26152;
              imag_value=19729;
            end
    4594  : begin
              real_value= 21600;
              imag_value=24630;
            end
    4595  : begin
              real_value= 16148;
              imag_value=28506;
            end
    4596  : begin
              real_value= 10021;
              imag_value=31191;
            end
    4597  : begin
              real_value= 3476;
              imag_value=32575;
            end
    4598  : begin
              real_value= -3210;
              imag_value=32603;
            end
    4599  : begin
              real_value= -9765;
              imag_value=31271;
            end
    4600  : begin
              real_value= -15914;
              imag_value=28636;
            end
    4601  : begin
              real_value= -21399;
              imag_value=24806;
            end
    4602  : begin
              real_value= -25990;
              imag_value=19943;
            end
    4603  : begin
              real_value= -29499;
              imag_value=14248;
            end
    4604  : begin
              real_value= -31779;
              imag_value=7959;
            end
    4605  : begin
              real_value= -32733;
              imag_value=1338;
            end
    4606  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    4607  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    4608  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    4609  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    4610  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    4611  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    4612  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    4613  : begin
              real_value= 802;
              imag_value=-32750;
            end
    4614  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    4615  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    4616  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    4617  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    4618  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    4619  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    4620  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    4621  : begin
              real_value= 32629;
              imag_value=2942;
            end
    4622  : begin
              real_value= 31351;
              imag_value=9508;
            end
    4623  : begin
              real_value= 28766;
              imag_value=15678;
            end
    4624  : begin
              real_value= 24981;
              imag_value=21194;
            end
    4625  : begin
              real_value= 20154;
              imag_value=25826;
            end
    4626  : begin
              real_value= 14489;
              imag_value=29382;
            end
    4627  : begin
              real_value= 8219;
              imag_value=31713;
            end
    4628  : begin
              real_value= 1606;
              imag_value=32721;
            end
    4629  : begin
              real_value= -5071;
              imag_value=32365;
            end
    4630  : begin
              real_value= -11539;
              imag_value=30661;
            end
    4631  : begin
              real_value= -17525;
              imag_value=27678;
            end
    4632  : begin
              real_value= -22782;
              imag_value=23541;
            end
    4633  : begin
              real_value= -27090;
              imag_value=18423;
            end
    4634  : begin
              real_value= -30267;
              imag_value=12537;
            end
    4635  : begin
              real_value= -32183;
              imag_value=6127;
            end
    4636  : begin
              real_value= -32757;
              imag_value=-535;
            end
    4637  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    4638  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    4639  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    4640  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    4641  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    4642  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    4643  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    4644  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    4645  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    4646  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    4647  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    4648  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    4649  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    4650  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    4651  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    4652  : begin
              real_value= 32407;
              imag_value=4806;
            end
    4653  : begin
              real_value= 30755;
              imag_value=11289;
            end
    4654  : begin
              real_value= 27820;
              imag_value=17299;
            end
    4655  : begin
              real_value= 23726;
              imag_value=22589;
            end
    4656  : begin
              real_value= 18644;
              imag_value=26938;
            end
    4657  : begin
              real_value= 12784;
              imag_value=30163;
            end
    4658  : begin
              real_value= 6390;
              imag_value=32131;
            end
    4659  : begin
              real_value= -267;
              imag_value=32759;
            end
    4660  : begin
              real_value= -6915;
              imag_value=32022;
            end
    4661  : begin
              real_value= -13274;
              imag_value=29950;
            end
    4662  : begin
              real_value= -19081;
              imag_value=26630;
            end
    4663  : begin
              real_value= -24092;
              imag_value=22199;
            end
    4664  : begin
              real_value= -28100;
              imag_value=16842;
            end
    4665  : begin
              real_value= -30935;
              imag_value=10783;
            end
    4666  : begin
              real_value= -32481;
              imag_value=4275;
            end
    4667  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    4668  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    4669  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    4670  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    4671  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    4672  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    4673  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    4674  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    4675  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    4676  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    4677  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    4678  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    4679  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    4680  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    4681  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    4682  : begin
              real_value= 32760;
              imag_value=0;
            end
    4683  : begin
              real_value= 32077;
              imag_value=6654;
            end
    4684  : begin
              real_value= 30057;
              imag_value=13030;
            end
    4685  : begin
              real_value= 26784;
              imag_value=18863;
            end
    4686  : begin
              real_value= 22395;
              imag_value=23911;
            end
    4687  : begin
              real_value= 17072;
              imag_value=27961;
            end
    4688  : begin
              real_value= 11036;
              imag_value=30846;
            end
    4689  : begin
              real_value= 4540;
              imag_value=32445;
            end
    4690  : begin
              real_value= -2142;
              imag_value=32691;
            end
    4691  : begin
              real_value= -8737;
              imag_value=31575;
            end
    4692  : begin
              real_value= -14968;
              imag_value=29142;
            end
    4693  : begin
              real_value= -20575;
              imag_value=25494;
            end
    4694  : begin
              real_value= -25324;
              imag_value=20783;
            end
    4695  : begin
              real_value= -29017;
              imag_value=15206;
            end
    4696  : begin
              real_value= -31501;
              imag_value=8995;
            end
    4697  : begin
              real_value= -32673;
              imag_value=2408;
            end
    4698  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    4699  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    4700  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    4701  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    4702  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    4703  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    4704  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    4705  : begin
              real_value= -267;
              imag_value=-32759;
            end
    4706  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    4707  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    4708  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    4709  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    4710  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    4711  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    4712  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    4713  : begin
              real_value= 32707;
              imag_value=1874;
            end
    4714  : begin
              real_value= 31645;
              imag_value=8477;
            end
    4715  : begin
              real_value= 29263;
              imag_value=14728;
            end
    4716  : begin
              real_value= 25661;
              imag_value=20365;
            end
    4717  : begin
              real_value= 20988;
              imag_value=25154;
            end
    4718  : begin
              real_value= 15442;
              imag_value=28892;
            end
    4719  : begin
              real_value= 9253;
              imag_value=31426;
            end
    4720  : begin
              real_value= 2676;
              imag_value=32651;
            end
    4721  : begin
              real_value= -4009;
              imag_value=32515;
            end
    4722  : begin
              real_value= -10529;
              imag_value=31023;
            end
    4723  : begin
              real_value= -16611;
              imag_value=28236;
            end
    4724  : begin
              real_value= -22001;
              imag_value=24274;
            end
    4725  : begin
              real_value= -26472;
              imag_value=19299;
            end
    4726  : begin
              real_value= -29841;
              imag_value=13520;
            end
    4727  : begin
              real_value= -31965;
              imag_value=7177;
            end
    4728  : begin
              real_value= -32757;
              imag_value=535;
            end
    4729  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    4730  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    4731  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    4732  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    4733  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    4734  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    4735  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    4736  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    4737  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    4738  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    4739  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    4740  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    4741  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    4742  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    4743  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    4744  : begin
              real_value= 32547;
              imag_value=3742;
            end
    4745  : begin
              real_value= 31107;
              imag_value=10275;
            end
    4746  : begin
              real_value= 28371;
              imag_value=16380;
            end
    4747  : begin
              real_value= 24453;
              imag_value=21801;
            end
    4748  : begin
              real_value= 19515;
              imag_value=26314;
            end
    4749  : begin
              real_value= 13764;
              imag_value=29729;
            end
    4750  : begin
              real_value= 7438;
              imag_value=31905;
            end
    4751  : begin
              real_value= 802;
              imag_value=32750;
            end
    4752  : begin
              real_value= -5864;
              imag_value=32231;
            end
    4753  : begin
              real_value= -12288;
              imag_value=30369;
            end
    4754  : begin
              real_value= -18200;
              imag_value=27240;
            end
    4755  : begin
              real_value= -23354;
              imag_value=22974;
            end
    4756  : begin
              real_value= -27534;
              imag_value=17752;
            end
    4757  : begin
              real_value= -30565;
              imag_value=11790;
            end
    4758  : begin
              real_value= -32323;
              imag_value=5336;
            end
    4759  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    4760  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    4761  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    4762  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    4763  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    4764  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    4765  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    4766  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    4767  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    4768  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    4769  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    4770  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    4771  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    4772  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    4773  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    4774  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    4775  : begin
              real_value= 32278;
              imag_value=5599;
            end
    4776  : begin
              real_value= 30468;
              imag_value=12039;
            end
    4777  : begin
              real_value= 27387;
              imag_value=17977;
            end
    4778  : begin
              real_value= 23165;
              imag_value=23165;
            end
    4779  : begin
              real_value= 17977;
              imag_value=27387;
            end
    4780  : begin
              real_value= 12039;
              imag_value=30468;
            end
    4781  : begin
              real_value= 5599;
              imag_value=32278;
            end
    4782  : begin
              real_value= -1070;
              imag_value=32743;
            end
    4783  : begin
              real_value= -7699;
              imag_value=31843;
            end
    4784  : begin
              real_value= -14006;
              imag_value=29615;
            end
    4785  : begin
              real_value= -19729;
              imag_value=26152;
            end
    4786  : begin
              real_value= -24630;
              imag_value=21600;
            end
    4787  : begin
              real_value= -28506;
              imag_value=16148;
            end
    4788  : begin
              real_value= -31191;
              imag_value=10021;
            end
    4789  : begin
              real_value= -32575;
              imag_value=3476;
            end
    4790  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    4791  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    4792  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    4793  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    4794  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    4795  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    4796  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    4797  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    4798  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    4799  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    4800  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    4801  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    4802  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    4803  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    4804  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    4805  : begin
              real_value= 32750;
              imag_value=802;
            end
    4806  : begin
              real_value= 31905;
              imag_value=7438;
            end
    4807  : begin
              real_value= 29729;
              imag_value=13764;
            end
    4808  : begin
              real_value= 26314;
              imag_value=19515;
            end
    4809  : begin
              real_value= 21801;
              imag_value=24453;
            end
    4810  : begin
              real_value= 16380;
              imag_value=28371;
            end
    4811  : begin
              real_value= 10275;
              imag_value=31107;
            end
    4812  : begin
              real_value= 3742;
              imag_value=32547;
            end
    4813  : begin
              real_value= -2942;
              imag_value=32629;
            end
    4814  : begin
              real_value= -9508;
              imag_value=31351;
            end
    4815  : begin
              real_value= -15678;
              imag_value=28766;
            end
    4816  : begin
              real_value= -21194;
              imag_value=24981;
            end
    4817  : begin
              real_value= -25826;
              imag_value=20154;
            end
    4818  : begin
              real_value= -29382;
              imag_value=14489;
            end
    4819  : begin
              real_value= -31713;
              imag_value=8219;
            end
    4820  : begin
              real_value= -32721;
              imag_value=1606;
            end
    4821  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    4822  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    4823  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    4824  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    4825  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    4826  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    4827  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    4828  : begin
              real_value= 535;
              imag_value=-32757;
            end
    4829  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    4830  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    4831  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    4832  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    4833  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    4834  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    4835  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    4836  : begin
              real_value= 32651;
              imag_value=2676;
            end
    4837  : begin
              real_value= 31426;
              imag_value=9253;
            end
    4838  : begin
              real_value= 28892;
              imag_value=15442;
            end
    4839  : begin
              real_value= 25154;
              imag_value=20988;
            end
    4840  : begin
              real_value= 20365;
              imag_value=25661;
            end
    4841  : begin
              real_value= 14728;
              imag_value=29263;
            end
    4842  : begin
              real_value= 8477;
              imag_value=31645;
            end
    4843  : begin
              real_value= 1874;
              imag_value=32707;
            end
    4844  : begin
              real_value= -4806;
              imag_value=32407;
            end
    4845  : begin
              real_value= -11289;
              imag_value=30755;
            end
    4846  : begin
              real_value= -17299;
              imag_value=27820;
            end
    4847  : begin
              real_value= -22589;
              imag_value=23726;
            end
    4848  : begin
              real_value= -26938;
              imag_value=18644;
            end
    4849  : begin
              real_value= -30163;
              imag_value=12784;
            end
    4850  : begin
              real_value= -32131;
              imag_value=6390;
            end
    4851  : begin
              real_value= -32759;
              imag_value=-267;
            end
    4852  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    4853  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    4854  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    4855  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    4856  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    4857  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    4858  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    4859  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    4860  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    4861  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    4862  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    4863  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    4864  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    4865  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    4866  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    4867  : begin
              real_value= 32445;
              imag_value=4540;
            end
    4868  : begin
              real_value= 30846;
              imag_value=11036;
            end
    4869  : begin
              real_value= 27961;
              imag_value=17072;
            end
    4870  : begin
              real_value= 23911;
              imag_value=22395;
            end
    4871  : begin
              real_value= 18863;
              imag_value=26784;
            end
    4872  : begin
              real_value= 13030;
              imag_value=30057;
            end
    4873  : begin
              real_value= 6654;
              imag_value=32077;
            end
    4874  : begin
              real_value= 0;
              imag_value=32760;
            end
    4875  : begin
              real_value= -6654;
              imag_value=32077;
            end
    4876  : begin
              real_value= -13030;
              imag_value=30057;
            end
    4877  : begin
              real_value= -18863;
              imag_value=26784;
            end
    4878  : begin
              real_value= -23911;
              imag_value=22395;
            end
    4879  : begin
              real_value= -27961;
              imag_value=17072;
            end
    4880  : begin
              real_value= -30846;
              imag_value=11036;
            end
    4881  : begin
              real_value= -32445;
              imag_value=4540;
            end
    4882  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    4883  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    4884  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    4885  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    4886  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    4887  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    4888  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    4889  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    4890  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    4891  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    4892  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    4893  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    4894  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    4895  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    4896  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    4897  : begin
              real_value= 32759;
              imag_value=-267;
            end
    4898  : begin
              real_value= 32131;
              imag_value=6390;
            end
    4899  : begin
              real_value= 30163;
              imag_value=12784;
            end
    4900  : begin
              real_value= 26938;
              imag_value=18644;
            end
    4901  : begin
              real_value= 22589;
              imag_value=23726;
            end
    4902  : begin
              real_value= 17299;
              imag_value=27820;
            end
    4903  : begin
              real_value= 11289;
              imag_value=30755;
            end
    4904  : begin
              real_value= 4806;
              imag_value=32407;
            end
    4905  : begin
              real_value= -1874;
              imag_value=32707;
            end
    4906  : begin
              real_value= -8477;
              imag_value=31645;
            end
    4907  : begin
              real_value= -14728;
              imag_value=29263;
            end
    4908  : begin
              real_value= -20365;
              imag_value=25661;
            end
    4909  : begin
              real_value= -25154;
              imag_value=20988;
            end
    4910  : begin
              real_value= -28892;
              imag_value=15442;
            end
    4911  : begin
              real_value= -31426;
              imag_value=9253;
            end
    4912  : begin
              real_value= -32651;
              imag_value=2676;
            end
    4913  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    4914  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    4915  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    4916  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    4917  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    4918  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    4919  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    4920  : begin
              real_value= -535;
              imag_value=-32757;
            end
    4921  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    4922  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    4923  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    4924  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    4925  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    4926  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    4927  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    4928  : begin
              real_value= 32721;
              imag_value=1606;
            end
    4929  : begin
              real_value= 31713;
              imag_value=8219;
            end
    4930  : begin
              real_value= 29382;
              imag_value=14489;
            end
    4931  : begin
              real_value= 25826;
              imag_value=20154;
            end
    4932  : begin
              real_value= 21194;
              imag_value=24981;
            end
    4933  : begin
              real_value= 15678;
              imag_value=28766;
            end
    4934  : begin
              real_value= 9508;
              imag_value=31351;
            end
    4935  : begin
              real_value= 2942;
              imag_value=32629;
            end
    4936  : begin
              real_value= -3742;
              imag_value=32547;
            end
    4937  : begin
              real_value= -10275;
              imag_value=31107;
            end
    4938  : begin
              real_value= -16380;
              imag_value=28371;
            end
    4939  : begin
              real_value= -21801;
              imag_value=24453;
            end
    4940  : begin
              real_value= -26314;
              imag_value=19515;
            end
    4941  : begin
              real_value= -29729;
              imag_value=13764;
            end
    4942  : begin
              real_value= -31905;
              imag_value=7438;
            end
    4943  : begin
              real_value= -32750;
              imag_value=802;
            end
    4944  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    4945  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    4946  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    4947  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    4948  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    4949  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    4950  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    4951  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    4952  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    4953  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    4954  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    4955  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    4956  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    4957  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    4958  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    4959  : begin
              real_value= 32575;
              imag_value=3476;
            end
    4960  : begin
              real_value= 31191;
              imag_value=10021;
            end
    4961  : begin
              real_value= 28506;
              imag_value=16148;
            end
    4962  : begin
              real_value= 24630;
              imag_value=21600;
            end
    4963  : begin
              real_value= 19729;
              imag_value=26152;
            end
    4964  : begin
              real_value= 14006;
              imag_value=29615;
            end
    4965  : begin
              real_value= 7699;
              imag_value=31843;
            end
    4966  : begin
              real_value= 1070;
              imag_value=32743;
            end
    4967  : begin
              real_value= -5599;
              imag_value=32278;
            end
    4968  : begin
              real_value= -12039;
              imag_value=30468;
            end
    4969  : begin
              real_value= -17977;
              imag_value=27387;
            end
    4970  : begin
              real_value= -23165;
              imag_value=23165;
            end
    4971  : begin
              real_value= -27387;
              imag_value=17977;
            end
    4972  : begin
              real_value= -30468;
              imag_value=12039;
            end
    4973  : begin
              real_value= -32278;
              imag_value=5599;
            end
    4974  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    4975  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    4976  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    4977  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    4978  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    4979  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    4980  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    4981  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    4982  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    4983  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    4984  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    4985  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    4986  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    4987  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    4988  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    4989  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    4990  : begin
              real_value= 32323;
              imag_value=5336;
            end
    4991  : begin
              real_value= 30565;
              imag_value=11790;
            end
    4992  : begin
              real_value= 27534;
              imag_value=17752;
            end
    4993  : begin
              real_value= 23354;
              imag_value=22974;
            end
    4994  : begin
              real_value= 18200;
              imag_value=27240;
            end
    4995  : begin
              real_value= 12288;
              imag_value=30369;
            end
    4996  : begin
              real_value= 5864;
              imag_value=32231;
            end
    4997  : begin
              real_value= -802;
              imag_value=32750;
            end
    4998  : begin
              real_value= -7438;
              imag_value=31905;
            end
    4999  : begin
              real_value= -13764;
              imag_value=29729;
            end
    5000  : begin
              real_value= -19515;
              imag_value=26314;
            end
    5001  : begin
              real_value= -24453;
              imag_value=21801;
            end
    5002  : begin
              real_value= -28371;
              imag_value=16380;
            end
    5003  : begin
              real_value= -31107;
              imag_value=10275;
            end
    5004  : begin
              real_value= -32547;
              imag_value=3742;
            end
    5005  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    5006  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    5007  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    5008  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    5009  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    5010  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    5011  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    5012  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    5013  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    5014  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    5015  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    5016  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    5017  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    5018  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    5019  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    5020  : begin
              real_value= 32757;
              imag_value=535;
            end
    5021  : begin
              real_value= 31965;
              imag_value=7177;
            end
    5022  : begin
              real_value= 29841;
              imag_value=13520;
            end
    5023  : begin
              real_value= 26472;
              imag_value=19299;
            end
    5024  : begin
              real_value= 22001;
              imag_value=24274;
            end
    5025  : begin
              real_value= 16611;
              imag_value=28236;
            end
    5026  : begin
              real_value= 10529;
              imag_value=31023;
            end
    5027  : begin
              real_value= 4009;
              imag_value=32515;
            end
    5028  : begin
              real_value= -2676;
              imag_value=32651;
            end
    5029  : begin
              real_value= -9253;
              imag_value=31426;
            end
    5030  : begin
              real_value= -15442;
              imag_value=28892;
            end
    5031  : begin
              real_value= -20988;
              imag_value=25154;
            end
    5032  : begin
              real_value= -25661;
              imag_value=20365;
            end
    5033  : begin
              real_value= -29263;
              imag_value=14728;
            end
    5034  : begin
              real_value= -31645;
              imag_value=8477;
            end
    5035  : begin
              real_value= -32707;
              imag_value=1874;
            end
    5036  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    5037  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    5038  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    5039  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    5040  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    5041  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    5042  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    5043  : begin
              real_value= 267;
              imag_value=-32759;
            end
    5044  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    5045  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    5046  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    5047  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    5048  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    5049  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    5050  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    5051  : begin
              real_value= 32673;
              imag_value=2408;
            end
    5052  : begin
              real_value= 31501;
              imag_value=8995;
            end
    5053  : begin
              real_value= 29017;
              imag_value=15206;
            end
    5054  : begin
              real_value= 25324;
              imag_value=20783;
            end
    5055  : begin
              real_value= 20575;
              imag_value=25494;
            end
    5056  : begin
              real_value= 14968;
              imag_value=29142;
            end
    5057  : begin
              real_value= 8737;
              imag_value=31575;
            end
    5058  : begin
              real_value= 2142;
              imag_value=32691;
            end
    5059  : begin
              real_value= -4540;
              imag_value=32445;
            end
    5060  : begin
              real_value= -11036;
              imag_value=30846;
            end
    5061  : begin
              real_value= -17072;
              imag_value=27961;
            end
    5062  : begin
              real_value= -22395;
              imag_value=23911;
            end
    5063  : begin
              real_value= -26784;
              imag_value=18863;
            end
    5064  : begin
              real_value= -30057;
              imag_value=13030;
            end
    5065  : begin
              real_value= -32077;
              imag_value=6654;
            end
    5066  : begin
              real_value= -32760;
              imag_value=0;
            end
    5067  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    5068  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    5069  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    5070  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    5071  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    5072  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    5073  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    5074  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    5075  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    5076  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    5077  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    5078  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    5079  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    5080  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    5081  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    5082  : begin
              real_value= 32481;
              imag_value=4275;
            end
    5083  : begin
              real_value= 30935;
              imag_value=10783;
            end
    5084  : begin
              real_value= 28100;
              imag_value=16842;
            end
    5085  : begin
              real_value= 24092;
              imag_value=22199;
            end
    5086  : begin
              real_value= 19081;
              imag_value=26630;
            end
    5087  : begin
              real_value= 13274;
              imag_value=29950;
            end
    5088  : begin
              real_value= 6915;
              imag_value=32022;
            end
    5089  : begin
              real_value= 267;
              imag_value=32759;
            end
    5090  : begin
              real_value= -6390;
              imag_value=32131;
            end
    5091  : begin
              real_value= -12784;
              imag_value=30163;
            end
    5092  : begin
              real_value= -18644;
              imag_value=26938;
            end
    5093  : begin
              real_value= -23726;
              imag_value=22589;
            end
    5094  : begin
              real_value= -27820;
              imag_value=17299;
            end
    5095  : begin
              real_value= -30755;
              imag_value=11289;
            end
    5096  : begin
              real_value= -32407;
              imag_value=4806;
            end
    5097  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    5098  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    5099  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    5100  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    5101  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    5102  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    5103  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    5104  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    5105  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    5106  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    5107  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    5108  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    5109  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    5110  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    5111  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    5112  : begin
              real_value= 32757;
              imag_value=-535;
            end
    5113  : begin
              real_value= 32183;
              imag_value=6127;
            end
    5114  : begin
              real_value= 30267;
              imag_value=12537;
            end
    5115  : begin
              real_value= 27090;
              imag_value=18423;
            end
    5116  : begin
              real_value= 22782;
              imag_value=23541;
            end
    5117  : begin
              real_value= 17525;
              imag_value=27678;
            end
    5118  : begin
              real_value= 11539;
              imag_value=30661;
            end
    5119  : begin
              real_value= 5071;
              imag_value=32365;
            end
    5120  : begin
              real_value= -1606;
              imag_value=32721;
            end
    5121  : begin
              real_value= -8219;
              imag_value=31713;
            end
    5122  : begin
              real_value= -14489;
              imag_value=29382;
            end
    5123  : begin
              real_value= -20154;
              imag_value=25826;
            end
    5124  : begin
              real_value= -24981;
              imag_value=21194;
            end
    5125  : begin
              real_value= -28766;
              imag_value=15678;
            end
    5126  : begin
              real_value= -31351;
              imag_value=9508;
            end
    5127  : begin
              real_value= -32629;
              imag_value=2942;
            end
    5128  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    5129  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    5130  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    5131  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    5132  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    5133  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    5134  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    5135  : begin
              real_value= -802;
              imag_value=-32750;
            end
    5136  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    5137  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    5138  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    5139  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    5140  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    5141  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    5142  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    5143  : begin
              real_value= 32733;
              imag_value=1338;
            end
    5144  : begin
              real_value= 31779;
              imag_value=7959;
            end
    5145  : begin
              real_value= 29499;
              imag_value=14248;
            end
    5146  : begin
              real_value= 25990;
              imag_value=19943;
            end
    5147  : begin
              real_value= 21399;
              imag_value=24806;
            end
    5148  : begin
              real_value= 15914;
              imag_value=28636;
            end
    5149  : begin
              real_value= 9765;
              imag_value=31271;
            end
    5150  : begin
              real_value= 3210;
              imag_value=32603;
            end
    5151  : begin
              real_value= -3476;
              imag_value=32575;
            end
    5152  : begin
              real_value= -10021;
              imag_value=31191;
            end
    5153  : begin
              real_value= -16148;
              imag_value=28506;
            end
    5154  : begin
              real_value= -21600;
              imag_value=24630;
            end
    5155  : begin
              real_value= -26152;
              imag_value=19729;
            end
    5156  : begin
              real_value= -29615;
              imag_value=14006;
            end
    5157  : begin
              real_value= -31843;
              imag_value=7699;
            end
    5158  : begin
              real_value= -32743;
              imag_value=1070;
            end
    5159  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    5160  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    5161  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    5162  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    5163  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    5164  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    5165  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    5166  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    5167  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    5168  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    5169  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    5170  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    5171  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    5172  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    5173  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    5174  : begin
              real_value= 32603;
              imag_value=3210;
            end
    5175  : begin
              real_value= 31271;
              imag_value=9765;
            end
    5176  : begin
              real_value= 28636;
              imag_value=15914;
            end
    5177  : begin
              real_value= 24806;
              imag_value=21399;
            end
    5178  : begin
              real_value= 19943;
              imag_value=25990;
            end
    5179  : begin
              real_value= 14248;
              imag_value=29499;
            end
    5180  : begin
              real_value= 7959;
              imag_value=31779;
            end
    5181  : begin
              real_value= 1338;
              imag_value=32733;
            end
    5182  : begin
              real_value= -5336;
              imag_value=32323;
            end
    5183  : begin
              real_value= -11790;
              imag_value=30565;
            end
    5184  : begin
              real_value= -17752;
              imag_value=27534;
            end
    5185  : begin
              real_value= -22974;
              imag_value=23354;
            end
    5186  : begin
              real_value= -27240;
              imag_value=18200;
            end
    5187  : begin
              real_value= -30369;
              imag_value=12288;
            end
    5188  : begin
              real_value= -32231;
              imag_value=5864;
            end
    5189  : begin
              real_value= -32750;
              imag_value=-802;
            end
    5190  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    5191  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    5192  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    5193  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    5194  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    5195  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    5196  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    5197  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    5198  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    5199  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    5200  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    5201  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    5202  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    5203  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    5204  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    5205  : begin
              real_value= 32365;
              imag_value=5071;
            end
    5206  : begin
              real_value= 30661;
              imag_value=11539;
            end
    5207  : begin
              real_value= 27678;
              imag_value=17525;
            end
    5208  : begin
              real_value= 23541;
              imag_value=22782;
            end
    5209  : begin
              real_value= 18423;
              imag_value=27090;
            end
    5210  : begin
              real_value= 12537;
              imag_value=30267;
            end
    5211  : begin
              real_value= 6127;
              imag_value=32183;
            end
    5212  : begin
              real_value= -535;
              imag_value=32757;
            end
    5213  : begin
              real_value= -7177;
              imag_value=31965;
            end
    5214  : begin
              real_value= -13520;
              imag_value=29841;
            end
    5215  : begin
              real_value= -19299;
              imag_value=26472;
            end
    5216  : begin
              real_value= -24274;
              imag_value=22001;
            end
    5217  : begin
              real_value= -28236;
              imag_value=16611;
            end
    5218  : begin
              real_value= -31023;
              imag_value=10529;
            end
    5219  : begin
              real_value= -32515;
              imag_value=4009;
            end
    5220  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    5221  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    5222  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    5223  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    5224  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    5225  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    5226  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    5227  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    5228  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    5229  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    5230  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    5231  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    5232  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    5233  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    5234  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    5235  : begin
              real_value= 32759;
              imag_value=267;
            end
    5236  : begin
              real_value= 32022;
              imag_value=6915;
            end
    5237  : begin
              real_value= 29950;
              imag_value=13274;
            end
    5238  : begin
              real_value= 26630;
              imag_value=19081;
            end
    5239  : begin
              real_value= 22199;
              imag_value=24092;
            end
    5240  : begin
              real_value= 16842;
              imag_value=28100;
            end
    5241  : begin
              real_value= 10783;
              imag_value=30935;
            end
    5242  : begin
              real_value= 4275;
              imag_value=32481;
            end
    5243  : begin
              real_value= -2408;
              imag_value=32673;
            end
    5244  : begin
              real_value= -8995;
              imag_value=31501;
            end
    5245  : begin
              real_value= -15206;
              imag_value=29017;
            end
    5246  : begin
              real_value= -20783;
              imag_value=25324;
            end
    5247  : begin
              real_value= -25494;
              imag_value=20575;
            end
    5248  : begin
              real_value= -29142;
              imag_value=14968;
            end
    5249  : begin
              real_value= -31575;
              imag_value=8737;
            end
    5250  : begin
              real_value= -32691;
              imag_value=2142;
            end
    5251  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    5252  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    5253  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    5254  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    5255  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    5256  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    5257  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    5258  : begin
              real_value= 0;
              imag_value=-32760;
            end
    5259  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    5260  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    5261  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    5262  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    5263  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    5264  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    5265  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    5266  : begin
              real_value= 32691;
              imag_value=2142;
            end
    5267  : begin
              real_value= 31575;
              imag_value=8737;
            end
    5268  : begin
              real_value= 29142;
              imag_value=14968;
            end
    5269  : begin
              real_value= 25494;
              imag_value=20575;
            end
    5270  : begin
              real_value= 20783;
              imag_value=25324;
            end
    5271  : begin
              real_value= 15206;
              imag_value=29017;
            end
    5272  : begin
              real_value= 8995;
              imag_value=31501;
            end
    5273  : begin
              real_value= 2408;
              imag_value=32673;
            end
    5274  : begin
              real_value= -4275;
              imag_value=32481;
            end
    5275  : begin
              real_value= -10783;
              imag_value=30935;
            end
    5276  : begin
              real_value= -16842;
              imag_value=28100;
            end
    5277  : begin
              real_value= -22199;
              imag_value=24092;
            end
    5278  : begin
              real_value= -26630;
              imag_value=19081;
            end
    5279  : begin
              real_value= -29950;
              imag_value=13274;
            end
    5280  : begin
              real_value= -32022;
              imag_value=6915;
            end
    5281  : begin
              real_value= -32759;
              imag_value=267;
            end
    5282  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    5283  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    5284  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    5285  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    5286  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    5287  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    5288  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    5289  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    5290  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    5291  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    5292  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    5293  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    5294  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    5295  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    5296  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    5297  : begin
              real_value= 32515;
              imag_value=4009;
            end
    5298  : begin
              real_value= 31023;
              imag_value=10529;
            end
    5299  : begin
              real_value= 28236;
              imag_value=16611;
            end
    5300  : begin
              real_value= 24274;
              imag_value=22001;
            end
    5301  : begin
              real_value= 19299;
              imag_value=26472;
            end
    5302  : begin
              real_value= 13520;
              imag_value=29841;
            end
    5303  : begin
              real_value= 7177;
              imag_value=31965;
            end
    5304  : begin
              real_value= 535;
              imag_value=32757;
            end
    5305  : begin
              real_value= -6127;
              imag_value=32183;
            end
    5306  : begin
              real_value= -12537;
              imag_value=30267;
            end
    5307  : begin
              real_value= -18423;
              imag_value=27090;
            end
    5308  : begin
              real_value= -23541;
              imag_value=22782;
            end
    5309  : begin
              real_value= -27678;
              imag_value=17525;
            end
    5310  : begin
              real_value= -30661;
              imag_value=11539;
            end
    5311  : begin
              real_value= -32365;
              imag_value=5071;
            end
    5312  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    5313  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    5314  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    5315  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    5316  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    5317  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    5318  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    5319  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    5320  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    5321  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    5322  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    5323  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    5324  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    5325  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    5326  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    5327  : begin
              real_value= 32750;
              imag_value=-802;
            end
    5328  : begin
              real_value= 32231;
              imag_value=5864;
            end
    5329  : begin
              real_value= 30369;
              imag_value=12288;
            end
    5330  : begin
              real_value= 27240;
              imag_value=18200;
            end
    5331  : begin
              real_value= 22974;
              imag_value=23354;
            end
    5332  : begin
              real_value= 17752;
              imag_value=27534;
            end
    5333  : begin
              real_value= 11790;
              imag_value=30565;
            end
    5334  : begin
              real_value= 5336;
              imag_value=32323;
            end
    5335  : begin
              real_value= -1338;
              imag_value=32733;
            end
    5336  : begin
              real_value= -7959;
              imag_value=31779;
            end
    5337  : begin
              real_value= -14248;
              imag_value=29499;
            end
    5338  : begin
              real_value= -19943;
              imag_value=25990;
            end
    5339  : begin
              real_value= -24806;
              imag_value=21399;
            end
    5340  : begin
              real_value= -28636;
              imag_value=15914;
            end
    5341  : begin
              real_value= -31271;
              imag_value=9765;
            end
    5342  : begin
              real_value= -32603;
              imag_value=3210;
            end
    5343  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    5344  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    5345  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    5346  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    5347  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    5348  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    5349  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    5350  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    5351  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    5352  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    5353  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    5354  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    5355  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    5356  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    5357  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    5358  : begin
              real_value= 32743;
              imag_value=1070;
            end
    5359  : begin
              real_value= 31843;
              imag_value=7699;
            end
    5360  : begin
              real_value= 29615;
              imag_value=14006;
            end
    5361  : begin
              real_value= 26152;
              imag_value=19729;
            end
    5362  : begin
              real_value= 21600;
              imag_value=24630;
            end
    5363  : begin
              real_value= 16148;
              imag_value=28506;
            end
    5364  : begin
              real_value= 10021;
              imag_value=31191;
            end
    5365  : begin
              real_value= 3476;
              imag_value=32575;
            end
    5366  : begin
              real_value= -3210;
              imag_value=32603;
            end
    5367  : begin
              real_value= -9765;
              imag_value=31271;
            end
    5368  : begin
              real_value= -15914;
              imag_value=28636;
            end
    5369  : begin
              real_value= -21399;
              imag_value=24806;
            end
    5370  : begin
              real_value= -25990;
              imag_value=19943;
            end
    5371  : begin
              real_value= -29499;
              imag_value=14248;
            end
    5372  : begin
              real_value= -31779;
              imag_value=7959;
            end
    5373  : begin
              real_value= -32733;
              imag_value=1338;
            end
    5374  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    5375  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    5376  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    5377  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    5378  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    5379  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    5380  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    5381  : begin
              real_value= 802;
              imag_value=-32750;
            end
    5382  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    5383  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    5384  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    5385  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    5386  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    5387  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    5388  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    5389  : begin
              real_value= 32629;
              imag_value=2942;
            end
    5390  : begin
              real_value= 31351;
              imag_value=9508;
            end
    5391  : begin
              real_value= 28766;
              imag_value=15678;
            end
    5392  : begin
              real_value= 24981;
              imag_value=21194;
            end
    5393  : begin
              real_value= 20154;
              imag_value=25826;
            end
    5394  : begin
              real_value= 14489;
              imag_value=29382;
            end
    5395  : begin
              real_value= 8219;
              imag_value=31713;
            end
    5396  : begin
              real_value= 1606;
              imag_value=32721;
            end
    5397  : begin
              real_value= -5071;
              imag_value=32365;
            end
    5398  : begin
              real_value= -11539;
              imag_value=30661;
            end
    5399  : begin
              real_value= -17525;
              imag_value=27678;
            end
    5400  : begin
              real_value= -22782;
              imag_value=23541;
            end
    5401  : begin
              real_value= -27090;
              imag_value=18423;
            end
    5402  : begin
              real_value= -30267;
              imag_value=12537;
            end
    5403  : begin
              real_value= -32183;
              imag_value=6127;
            end
    5404  : begin
              real_value= -32757;
              imag_value=-535;
            end
    5405  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    5406  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    5407  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    5408  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    5409  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    5410  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    5411  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    5412  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    5413  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    5414  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    5415  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    5416  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    5417  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    5418  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    5419  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    5420  : begin
              real_value= 32407;
              imag_value=4806;
            end
    5421  : begin
              real_value= 30755;
              imag_value=11289;
            end
    5422  : begin
              real_value= 27820;
              imag_value=17299;
            end
    5423  : begin
              real_value= 23726;
              imag_value=22589;
            end
    5424  : begin
              real_value= 18644;
              imag_value=26938;
            end
    5425  : begin
              real_value= 12784;
              imag_value=30163;
            end
    5426  : begin
              real_value= 6390;
              imag_value=32131;
            end
    5427  : begin
              real_value= -267;
              imag_value=32759;
            end
    5428  : begin
              real_value= -6915;
              imag_value=32022;
            end
    5429  : begin
              real_value= -13274;
              imag_value=29950;
            end
    5430  : begin
              real_value= -19081;
              imag_value=26630;
            end
    5431  : begin
              real_value= -24092;
              imag_value=22199;
            end
    5432  : begin
              real_value= -28100;
              imag_value=16842;
            end
    5433  : begin
              real_value= -30935;
              imag_value=10783;
            end
    5434  : begin
              real_value= -32481;
              imag_value=4275;
            end
    5435  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    5436  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    5437  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    5438  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    5439  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    5440  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    5441  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    5442  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    5443  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    5444  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    5445  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    5446  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    5447  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    5448  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    5449  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    5450  : begin
              real_value= 32760;
              imag_value=0;
            end
    5451  : begin
              real_value= 32077;
              imag_value=6654;
            end
    5452  : begin
              real_value= 30057;
              imag_value=13030;
            end
    5453  : begin
              real_value= 26784;
              imag_value=18863;
            end
    5454  : begin
              real_value= 22395;
              imag_value=23911;
            end
    5455  : begin
              real_value= 17072;
              imag_value=27961;
            end
    5456  : begin
              real_value= 11036;
              imag_value=30846;
            end
    5457  : begin
              real_value= 4540;
              imag_value=32445;
            end
    5458  : begin
              real_value= -2142;
              imag_value=32691;
            end
    5459  : begin
              real_value= -8737;
              imag_value=31575;
            end
    5460  : begin
              real_value= -14968;
              imag_value=29142;
            end
    5461  : begin
              real_value= -20575;
              imag_value=25494;
            end
    5462  : begin
              real_value= -25324;
              imag_value=20783;
            end
    5463  : begin
              real_value= -29017;
              imag_value=15206;
            end
    5464  : begin
              real_value= -31501;
              imag_value=8995;
            end
    5465  : begin
              real_value= -32673;
              imag_value=2408;
            end
    5466  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    5467  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    5468  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    5469  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    5470  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    5471  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    5472  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    5473  : begin
              real_value= -267;
              imag_value=-32759;
            end
    5474  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    5475  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    5476  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    5477  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    5478  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    5479  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    5480  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    5481  : begin
              real_value= 32707;
              imag_value=1874;
            end
    5482  : begin
              real_value= 31645;
              imag_value=8477;
            end
    5483  : begin
              real_value= 29263;
              imag_value=14728;
            end
    5484  : begin
              real_value= 25661;
              imag_value=20365;
            end
    5485  : begin
              real_value= 20988;
              imag_value=25154;
            end
    5486  : begin
              real_value= 15442;
              imag_value=28892;
            end
    5487  : begin
              real_value= 9253;
              imag_value=31426;
            end
    5488  : begin
              real_value= 2676;
              imag_value=32651;
            end
    5489  : begin
              real_value= -4009;
              imag_value=32515;
            end
    5490  : begin
              real_value= -10529;
              imag_value=31023;
            end
    5491  : begin
              real_value= -16611;
              imag_value=28236;
            end
    5492  : begin
              real_value= -22001;
              imag_value=24274;
            end
    5493  : begin
              real_value= -26472;
              imag_value=19299;
            end
    5494  : begin
              real_value= -29841;
              imag_value=13520;
            end
    5495  : begin
              real_value= -31965;
              imag_value=7177;
            end
    5496  : begin
              real_value= -32757;
              imag_value=535;
            end
    5497  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    5498  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    5499  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    5500  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    5501  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    5502  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    5503  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    5504  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    5505  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    5506  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    5507  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    5508  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    5509  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    5510  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    5511  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    5512  : begin
              real_value= 32547;
              imag_value=3742;
            end
    5513  : begin
              real_value= 31107;
              imag_value=10275;
            end
    5514  : begin
              real_value= 28371;
              imag_value=16380;
            end
    5515  : begin
              real_value= 24453;
              imag_value=21801;
            end
    5516  : begin
              real_value= 19515;
              imag_value=26314;
            end
    5517  : begin
              real_value= 13764;
              imag_value=29729;
            end
    5518  : begin
              real_value= 7438;
              imag_value=31905;
            end
    5519  : begin
              real_value= 802;
              imag_value=32750;
            end
    5520  : begin
              real_value= -5864;
              imag_value=32231;
            end
    5521  : begin
              real_value= -12288;
              imag_value=30369;
            end
    5522  : begin
              real_value= -18200;
              imag_value=27240;
            end
    5523  : begin
              real_value= -23354;
              imag_value=22974;
            end
    5524  : begin
              real_value= -27534;
              imag_value=17752;
            end
    5525  : begin
              real_value= -30565;
              imag_value=11790;
            end
    5526  : begin
              real_value= -32323;
              imag_value=5336;
            end
    5527  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    5528  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    5529  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    5530  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    5531  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    5532  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    5533  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    5534  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    5535  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    5536  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    5537  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    5538  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    5539  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    5540  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    5541  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    5542  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    5543  : begin
              real_value= 32278;
              imag_value=5599;
            end
    5544  : begin
              real_value= 30468;
              imag_value=12039;
            end
    5545  : begin
              real_value= 27387;
              imag_value=17977;
            end
    5546  : begin
              real_value= 23165;
              imag_value=23165;
            end
    5547  : begin
              real_value= 17977;
              imag_value=27387;
            end
    5548  : begin
              real_value= 12039;
              imag_value=30468;
            end
    5549  : begin
              real_value= 5599;
              imag_value=32278;
            end
    5550  : begin
              real_value= -1070;
              imag_value=32743;
            end
    5551  : begin
              real_value= -7699;
              imag_value=31843;
            end
    5552  : begin
              real_value= -14006;
              imag_value=29615;
            end
    5553  : begin
              real_value= -19729;
              imag_value=26152;
            end
    5554  : begin
              real_value= -24630;
              imag_value=21600;
            end
    5555  : begin
              real_value= -28506;
              imag_value=16148;
            end
    5556  : begin
              real_value= -31191;
              imag_value=10021;
            end
    5557  : begin
              real_value= -32575;
              imag_value=3476;
            end
    5558  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    5559  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    5560  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    5561  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    5562  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    5563  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    5564  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    5565  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    5566  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    5567  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    5568  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    5569  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    5570  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    5571  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    5572  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    5573  : begin
              real_value= 32750;
              imag_value=802;
            end
    5574  : begin
              real_value= 31905;
              imag_value=7438;
            end
    5575  : begin
              real_value= 29729;
              imag_value=13764;
            end
    5576  : begin
              real_value= 26314;
              imag_value=19515;
            end
    5577  : begin
              real_value= 21801;
              imag_value=24453;
            end
    5578  : begin
              real_value= 16380;
              imag_value=28371;
            end
    5579  : begin
              real_value= 10275;
              imag_value=31107;
            end
    5580  : begin
              real_value= 3742;
              imag_value=32547;
            end
    5581  : begin
              real_value= -2942;
              imag_value=32629;
            end
    5582  : begin
              real_value= -9508;
              imag_value=31351;
            end
    5583  : begin
              real_value= -15678;
              imag_value=28766;
            end
    5584  : begin
              real_value= -21194;
              imag_value=24981;
            end
    5585  : begin
              real_value= -25826;
              imag_value=20154;
            end
    5586  : begin
              real_value= -29382;
              imag_value=14489;
            end
    5587  : begin
              real_value= -31713;
              imag_value=8219;
            end
    5588  : begin
              real_value= -32721;
              imag_value=1606;
            end
    5589  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    5590  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    5591  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    5592  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    5593  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    5594  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    5595  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    5596  : begin
              real_value= 535;
              imag_value=-32757;
            end
    5597  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    5598  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    5599  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    5600  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    5601  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    5602  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    5603  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    5604  : begin
              real_value= 32651;
              imag_value=2676;
            end
    5605  : begin
              real_value= 31426;
              imag_value=9253;
            end
    5606  : begin
              real_value= 28892;
              imag_value=15442;
            end
    5607  : begin
              real_value= 25154;
              imag_value=20988;
            end
    5608  : begin
              real_value= 20365;
              imag_value=25661;
            end
    5609  : begin
              real_value= 14728;
              imag_value=29263;
            end
    5610  : begin
              real_value= 8477;
              imag_value=31645;
            end
    5611  : begin
              real_value= 1874;
              imag_value=32707;
            end
    5612  : begin
              real_value= -4806;
              imag_value=32407;
            end
    5613  : begin
              real_value= -11289;
              imag_value=30755;
            end
    5614  : begin
              real_value= -17299;
              imag_value=27820;
            end
    5615  : begin
              real_value= -22589;
              imag_value=23726;
            end
    5616  : begin
              real_value= -26938;
              imag_value=18644;
            end
    5617  : begin
              real_value= -30163;
              imag_value=12784;
            end
    5618  : begin
              real_value= -32131;
              imag_value=6390;
            end
    5619  : begin
              real_value= -32759;
              imag_value=-267;
            end
    5620  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    5621  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    5622  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    5623  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    5624  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    5625  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    5626  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    5627  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    5628  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    5629  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    5630  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    5631  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    5632  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    5633  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    5634  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    5635  : begin
              real_value= 32445;
              imag_value=4540;
            end
    5636  : begin
              real_value= 30846;
              imag_value=11036;
            end
    5637  : begin
              real_value= 27961;
              imag_value=17072;
            end
    5638  : begin
              real_value= 23911;
              imag_value=22395;
            end
    5639  : begin
              real_value= 18863;
              imag_value=26784;
            end
    5640  : begin
              real_value= 13030;
              imag_value=30057;
            end
    5641  : begin
              real_value= 6654;
              imag_value=32077;
            end
    5642  : begin
              real_value= 0;
              imag_value=32760;
            end
    5643  : begin
              real_value= -6654;
              imag_value=32077;
            end
    5644  : begin
              real_value= -13030;
              imag_value=30057;
            end
    5645  : begin
              real_value= -18863;
              imag_value=26784;
            end
    5646  : begin
              real_value= -23911;
              imag_value=22395;
            end
    5647  : begin
              real_value= -27961;
              imag_value=17072;
            end
    5648  : begin
              real_value= -30846;
              imag_value=11036;
            end
    5649  : begin
              real_value= -32445;
              imag_value=4540;
            end
    5650  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    5651  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    5652  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    5653  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    5654  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    5655  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    5656  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    5657  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    5658  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    5659  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    5660  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    5661  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    5662  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    5663  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    5664  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    5665  : begin
              real_value= 32759;
              imag_value=-267;
            end
    5666  : begin
              real_value= 32131;
              imag_value=6390;
            end
    5667  : begin
              real_value= 30163;
              imag_value=12784;
            end
    5668  : begin
              real_value= 26938;
              imag_value=18644;
            end
    5669  : begin
              real_value= 22589;
              imag_value=23726;
            end
    5670  : begin
              real_value= 17299;
              imag_value=27820;
            end
    5671  : begin
              real_value= 11289;
              imag_value=30755;
            end
    5672  : begin
              real_value= 4806;
              imag_value=32407;
            end
    5673  : begin
              real_value= -1874;
              imag_value=32707;
            end
    5674  : begin
              real_value= -8477;
              imag_value=31645;
            end
    5675  : begin
              real_value= -14728;
              imag_value=29263;
            end
    5676  : begin
              real_value= -20365;
              imag_value=25661;
            end
    5677  : begin
              real_value= -25154;
              imag_value=20988;
            end
    5678  : begin
              real_value= -28892;
              imag_value=15442;
            end
    5679  : begin
              real_value= -31426;
              imag_value=9253;
            end
    5680  : begin
              real_value= -32651;
              imag_value=2676;
            end
    5681  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    5682  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    5683  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    5684  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    5685  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    5686  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    5687  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    5688  : begin
              real_value= -535;
              imag_value=-32757;
            end
    5689  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    5690  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    5691  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    5692  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    5693  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    5694  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    5695  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    5696  : begin
              real_value= 32721;
              imag_value=1606;
            end
    5697  : begin
              real_value= 31713;
              imag_value=8219;
            end
    5698  : begin
              real_value= 29382;
              imag_value=14489;
            end
    5699  : begin
              real_value= 25826;
              imag_value=20154;
            end
    5700  : begin
              real_value= 21194;
              imag_value=24981;
            end
    5701  : begin
              real_value= 15678;
              imag_value=28766;
            end
    5702  : begin
              real_value= 9508;
              imag_value=31351;
            end
    5703  : begin
              real_value= 2942;
              imag_value=32629;
            end
    5704  : begin
              real_value= -3742;
              imag_value=32547;
            end
    5705  : begin
              real_value= -10275;
              imag_value=31107;
            end
    5706  : begin
              real_value= -16380;
              imag_value=28371;
            end
    5707  : begin
              real_value= -21801;
              imag_value=24453;
            end
    5708  : begin
              real_value= -26314;
              imag_value=19515;
            end
    5709  : begin
              real_value= -29729;
              imag_value=13764;
            end
    5710  : begin
              real_value= -31905;
              imag_value=7438;
            end
    5711  : begin
              real_value= -32750;
              imag_value=802;
            end
    5712  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    5713  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    5714  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    5715  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    5716  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    5717  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    5718  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    5719  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    5720  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    5721  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    5722  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    5723  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    5724  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    5725  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    5726  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    5727  : begin
              real_value= 32575;
              imag_value=3476;
            end
    5728  : begin
              real_value= 31191;
              imag_value=10021;
            end
    5729  : begin
              real_value= 28506;
              imag_value=16148;
            end
    5730  : begin
              real_value= 24630;
              imag_value=21600;
            end
    5731  : begin
              real_value= 19729;
              imag_value=26152;
            end
    5732  : begin
              real_value= 14006;
              imag_value=29615;
            end
    5733  : begin
              real_value= 7699;
              imag_value=31843;
            end
    5734  : begin
              real_value= 1070;
              imag_value=32743;
            end
    5735  : begin
              real_value= -5599;
              imag_value=32278;
            end
    5736  : begin
              real_value= -12039;
              imag_value=30468;
            end
    5737  : begin
              real_value= -17977;
              imag_value=27387;
            end
    5738  : begin
              real_value= -23165;
              imag_value=23165;
            end
    5739  : begin
              real_value= -27387;
              imag_value=17977;
            end
    5740  : begin
              real_value= -30468;
              imag_value=12039;
            end
    5741  : begin
              real_value= -32278;
              imag_value=5599;
            end
    5742  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    5743  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    5744  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    5745  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    5746  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    5747  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    5748  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    5749  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    5750  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    5751  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    5752  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    5753  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    5754  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    5755  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    5756  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    5757  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    5758  : begin
              real_value= 32323;
              imag_value=5336;
            end
    5759  : begin
              real_value= 30565;
              imag_value=11790;
            end
    5760  : begin
              real_value= 27534;
              imag_value=17752;
            end
    5761  : begin
              real_value= 23354;
              imag_value=22974;
            end
    5762  : begin
              real_value= 18200;
              imag_value=27240;
            end
    5763  : begin
              real_value= 12288;
              imag_value=30369;
            end
    5764  : begin
              real_value= 5864;
              imag_value=32231;
            end
    5765  : begin
              real_value= -802;
              imag_value=32750;
            end
    5766  : begin
              real_value= -7438;
              imag_value=31905;
            end
    5767  : begin
              real_value= -13764;
              imag_value=29729;
            end
    5768  : begin
              real_value= -19515;
              imag_value=26314;
            end
    5769  : begin
              real_value= -24453;
              imag_value=21801;
            end
    5770  : begin
              real_value= -28371;
              imag_value=16380;
            end
    5771  : begin
              real_value= -31107;
              imag_value=10275;
            end
    5772  : begin
              real_value= -32547;
              imag_value=3742;
            end
    5773  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    5774  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    5775  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    5776  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    5777  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    5778  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    5779  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    5780  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    5781  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    5782  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    5783  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    5784  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    5785  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    5786  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    5787  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    5788  : begin
              real_value= 32757;
              imag_value=535;
            end
    5789  : begin
              real_value= 31965;
              imag_value=7177;
            end
    5790  : begin
              real_value= 29841;
              imag_value=13520;
            end
    5791  : begin
              real_value= 26472;
              imag_value=19299;
            end
    5792  : begin
              real_value= 22001;
              imag_value=24274;
            end
    5793  : begin
              real_value= 16611;
              imag_value=28236;
            end
    5794  : begin
              real_value= 10529;
              imag_value=31023;
            end
    5795  : begin
              real_value= 4009;
              imag_value=32515;
            end
    5796  : begin
              real_value= -2676;
              imag_value=32651;
            end
    5797  : begin
              real_value= -9253;
              imag_value=31426;
            end
    5798  : begin
              real_value= -15442;
              imag_value=28892;
            end
    5799  : begin
              real_value= -20988;
              imag_value=25154;
            end
    5800  : begin
              real_value= -25661;
              imag_value=20365;
            end
    5801  : begin
              real_value= -29263;
              imag_value=14728;
            end
    5802  : begin
              real_value= -31645;
              imag_value=8477;
            end
    5803  : begin
              real_value= -32707;
              imag_value=1874;
            end
    5804  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    5805  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    5806  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    5807  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    5808  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    5809  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    5810  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    5811  : begin
              real_value= 267;
              imag_value=-32759;
            end
    5812  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    5813  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    5814  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    5815  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    5816  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    5817  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    5818  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    5819  : begin
              real_value= 32673;
              imag_value=2408;
            end
    5820  : begin
              real_value= 31501;
              imag_value=8995;
            end
    5821  : begin
              real_value= 29017;
              imag_value=15206;
            end
    5822  : begin
              real_value= 25324;
              imag_value=20783;
            end
    5823  : begin
              real_value= 20575;
              imag_value=25494;
            end
    5824  : begin
              real_value= 14968;
              imag_value=29142;
            end
    5825  : begin
              real_value= 8737;
              imag_value=31575;
            end
    5826  : begin
              real_value= 2142;
              imag_value=32691;
            end
    5827  : begin
              real_value= -4540;
              imag_value=32445;
            end
    5828  : begin
              real_value= -11036;
              imag_value=30846;
            end
    5829  : begin
              real_value= -17072;
              imag_value=27961;
            end
    5830  : begin
              real_value= -22395;
              imag_value=23911;
            end
    5831  : begin
              real_value= -26784;
              imag_value=18863;
            end
    5832  : begin
              real_value= -30057;
              imag_value=13030;
            end
    5833  : begin
              real_value= -32077;
              imag_value=6654;
            end
    5834  : begin
              real_value= -32760;
              imag_value=0;
            end
    5835  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    5836  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    5837  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    5838  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    5839  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    5840  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    5841  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    5842  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    5843  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    5844  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    5845  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    5846  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    5847  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    5848  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    5849  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    5850  : begin
              real_value= 32481;
              imag_value=4275;
            end
    5851  : begin
              real_value= 30935;
              imag_value=10783;
            end
    5852  : begin
              real_value= 28100;
              imag_value=16842;
            end
    5853  : begin
              real_value= 24092;
              imag_value=22199;
            end
    5854  : begin
              real_value= 19081;
              imag_value=26630;
            end
    5855  : begin
              real_value= 13274;
              imag_value=29950;
            end
    5856  : begin
              real_value= 6915;
              imag_value=32022;
            end
    5857  : begin
              real_value= 267;
              imag_value=32759;
            end
    5858  : begin
              real_value= -6390;
              imag_value=32131;
            end
    5859  : begin
              real_value= -12784;
              imag_value=30163;
            end
    5860  : begin
              real_value= -18644;
              imag_value=26938;
            end
    5861  : begin
              real_value= -23726;
              imag_value=22589;
            end
    5862  : begin
              real_value= -27820;
              imag_value=17299;
            end
    5863  : begin
              real_value= -30755;
              imag_value=11289;
            end
    5864  : begin
              real_value= -32407;
              imag_value=4806;
            end
    5865  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    5866  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    5867  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    5868  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    5869  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    5870  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    5871  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    5872  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    5873  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    5874  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    5875  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    5876  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    5877  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    5878  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    5879  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    5880  : begin
              real_value= 32757;
              imag_value=-535;
            end
    5881  : begin
              real_value= 32183;
              imag_value=6127;
            end
    5882  : begin
              real_value= 30267;
              imag_value=12537;
            end
    5883  : begin
              real_value= 27090;
              imag_value=18423;
            end
    5884  : begin
              real_value= 22782;
              imag_value=23541;
            end
    5885  : begin
              real_value= 17525;
              imag_value=27678;
            end
    5886  : begin
              real_value= 11539;
              imag_value=30661;
            end
    5887  : begin
              real_value= 5071;
              imag_value=32365;
            end
    5888  : begin
              real_value= -1606;
              imag_value=32721;
            end
    5889  : begin
              real_value= -8219;
              imag_value=31713;
            end
    5890  : begin
              real_value= -14489;
              imag_value=29382;
            end
    5891  : begin
              real_value= -20154;
              imag_value=25826;
            end
    5892  : begin
              real_value= -24981;
              imag_value=21194;
            end
    5893  : begin
              real_value= -28766;
              imag_value=15678;
            end
    5894  : begin
              real_value= -31351;
              imag_value=9508;
            end
    5895  : begin
              real_value= -32629;
              imag_value=2942;
            end
    5896  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    5897  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    5898  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    5899  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    5900  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    5901  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    5902  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    5903  : begin
              real_value= -802;
              imag_value=-32750;
            end
    5904  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    5905  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    5906  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    5907  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    5908  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    5909  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    5910  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    5911  : begin
              real_value= 32733;
              imag_value=1338;
            end
    5912  : begin
              real_value= 31779;
              imag_value=7959;
            end
    5913  : begin
              real_value= 29499;
              imag_value=14248;
            end
    5914  : begin
              real_value= 25990;
              imag_value=19943;
            end
    5915  : begin
              real_value= 21399;
              imag_value=24806;
            end
    5916  : begin
              real_value= 15914;
              imag_value=28636;
            end
    5917  : begin
              real_value= 9765;
              imag_value=31271;
            end
    5918  : begin
              real_value= 3210;
              imag_value=32603;
            end
    5919  : begin
              real_value= -3476;
              imag_value=32575;
            end
    5920  : begin
              real_value= -10021;
              imag_value=31191;
            end
    5921  : begin
              real_value= -16148;
              imag_value=28506;
            end
    5922  : begin
              real_value= -21600;
              imag_value=24630;
            end
    5923  : begin
              real_value= -26152;
              imag_value=19729;
            end
    5924  : begin
              real_value= -29615;
              imag_value=14006;
            end
    5925  : begin
              real_value= -31843;
              imag_value=7699;
            end
    5926  : begin
              real_value= -32743;
              imag_value=1070;
            end
    5927  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    5928  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    5929  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    5930  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    5931  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    5932  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    5933  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    5934  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    5935  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    5936  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    5937  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    5938  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    5939  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    5940  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    5941  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    5942  : begin
              real_value= 32603;
              imag_value=3210;
            end
    5943  : begin
              real_value= 31271;
              imag_value=9765;
            end
    5944  : begin
              real_value= 28636;
              imag_value=15914;
            end
    5945  : begin
              real_value= 24806;
              imag_value=21399;
            end
    5946  : begin
              real_value= 19943;
              imag_value=25990;
            end
    5947  : begin
              real_value= 14248;
              imag_value=29499;
            end
    5948  : begin
              real_value= 7959;
              imag_value=31779;
            end
    5949  : begin
              real_value= 1338;
              imag_value=32733;
            end
    5950  : begin
              real_value= -5336;
              imag_value=32323;
            end
    5951  : begin
              real_value= -11790;
              imag_value=30565;
            end
    5952  : begin
              real_value= -17752;
              imag_value=27534;
            end
    5953  : begin
              real_value= -22974;
              imag_value=23354;
            end
    5954  : begin
              real_value= -27240;
              imag_value=18200;
            end
    5955  : begin
              real_value= -30369;
              imag_value=12288;
            end
    5956  : begin
              real_value= -32231;
              imag_value=5864;
            end
    5957  : begin
              real_value= -32750;
              imag_value=-802;
            end
    5958  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    5959  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    5960  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    5961  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    5962  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    5963  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    5964  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    5965  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    5966  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    5967  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    5968  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    5969  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    5970  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    5971  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    5972  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    5973  : begin
              real_value= 32365;
              imag_value=5071;
            end
    5974  : begin
              real_value= 30661;
              imag_value=11539;
            end
    5975  : begin
              real_value= 27678;
              imag_value=17525;
            end
    5976  : begin
              real_value= 23541;
              imag_value=22782;
            end
    5977  : begin
              real_value= 18423;
              imag_value=27090;
            end
    5978  : begin
              real_value= 12537;
              imag_value=30267;
            end
    5979  : begin
              real_value= 6127;
              imag_value=32183;
            end
    5980  : begin
              real_value= -535;
              imag_value=32757;
            end
    5981  : begin
              real_value= -7177;
              imag_value=31965;
            end
    5982  : begin
              real_value= -13520;
              imag_value=29841;
            end
    5983  : begin
              real_value= -19299;
              imag_value=26472;
            end
    5984  : begin
              real_value= -24274;
              imag_value=22001;
            end
    5985  : begin
              real_value= -28236;
              imag_value=16611;
            end
    5986  : begin
              real_value= -31023;
              imag_value=10529;
            end
    5987  : begin
              real_value= -32515;
              imag_value=4009;
            end
    5988  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    5989  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    5990  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    5991  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    5992  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    5993  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    5994  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    5995  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    5996  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    5997  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    5998  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    5999  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    6000  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    6001  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    6002  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    6003  : begin
              real_value= 32759;
              imag_value=267;
            end
    6004  : begin
              real_value= 32022;
              imag_value=6915;
            end
    6005  : begin
              real_value= 29950;
              imag_value=13274;
            end
    6006  : begin
              real_value= 26630;
              imag_value=19081;
            end
    6007  : begin
              real_value= 22199;
              imag_value=24092;
            end
    6008  : begin
              real_value= 16842;
              imag_value=28100;
            end
    6009  : begin
              real_value= 10783;
              imag_value=30935;
            end
    6010  : begin
              real_value= 4275;
              imag_value=32481;
            end
    6011  : begin
              real_value= -2408;
              imag_value=32673;
            end
    6012  : begin
              real_value= -8995;
              imag_value=31501;
            end
    6013  : begin
              real_value= -15206;
              imag_value=29017;
            end
    6014  : begin
              real_value= -20783;
              imag_value=25324;
            end
    6015  : begin
              real_value= -25494;
              imag_value=20575;
            end
    6016  : begin
              real_value= -29142;
              imag_value=14968;
            end
    6017  : begin
              real_value= -31575;
              imag_value=8737;
            end
    6018  : begin
              real_value= -32691;
              imag_value=2142;
            end
    6019  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    6020  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    6021  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    6022  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    6023  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    6024  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    6025  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    6026  : begin
              real_value= 0;
              imag_value=-32760;
            end
    6027  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    6028  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    6029  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    6030  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    6031  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    6032  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    6033  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    6034  : begin
              real_value= 32691;
              imag_value=2142;
            end
    6035  : begin
              real_value= 31575;
              imag_value=8737;
            end
    6036  : begin
              real_value= 29142;
              imag_value=14968;
            end
    6037  : begin
              real_value= 25494;
              imag_value=20575;
            end
    6038  : begin
              real_value= 20783;
              imag_value=25324;
            end
    6039  : begin
              real_value= 15206;
              imag_value=29017;
            end
    6040  : begin
              real_value= 8995;
              imag_value=31501;
            end
    6041  : begin
              real_value= 2408;
              imag_value=32673;
            end
    6042  : begin
              real_value= -4275;
              imag_value=32481;
            end
    6043  : begin
              real_value= -10783;
              imag_value=30935;
            end
    6044  : begin
              real_value= -16842;
              imag_value=28100;
            end
    6045  : begin
              real_value= -22199;
              imag_value=24092;
            end
    6046  : begin
              real_value= -26630;
              imag_value=19081;
            end
    6047  : begin
              real_value= -29950;
              imag_value=13274;
            end
    6048  : begin
              real_value= -32022;
              imag_value=6915;
            end
    6049  : begin
              real_value= -32759;
              imag_value=267;
            end
    6050  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    6051  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    6052  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    6053  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    6054  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    6055  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    6056  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    6057  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    6058  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    6059  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    6060  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    6061  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    6062  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    6063  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    6064  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    6065  : begin
              real_value= 32515;
              imag_value=4009;
            end
    6066  : begin
              real_value= 31023;
              imag_value=10529;
            end
    6067  : begin
              real_value= 28236;
              imag_value=16611;
            end
    6068  : begin
              real_value= 24274;
              imag_value=22001;
            end
    6069  : begin
              real_value= 19299;
              imag_value=26472;
            end
    6070  : begin
              real_value= 13520;
              imag_value=29841;
            end
    6071  : begin
              real_value= 7177;
              imag_value=31965;
            end
    6072  : begin
              real_value= 535;
              imag_value=32757;
            end
    6073  : begin
              real_value= -6127;
              imag_value=32183;
            end
    6074  : begin
              real_value= -12537;
              imag_value=30267;
            end
    6075  : begin
              real_value= -18423;
              imag_value=27090;
            end
    6076  : begin
              real_value= -23541;
              imag_value=22782;
            end
    6077  : begin
              real_value= -27678;
              imag_value=17525;
            end
    6078  : begin
              real_value= -30661;
              imag_value=11539;
            end
    6079  : begin
              real_value= -32365;
              imag_value=5071;
            end
    6080  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    6081  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    6082  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    6083  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    6084  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    6085  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    6086  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    6087  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    6088  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    6089  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    6090  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    6091  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    6092  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    6093  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    6094  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    6095  : begin
              real_value= 32750;
              imag_value=-802;
            end
    6096  : begin
              real_value= 32231;
              imag_value=5864;
            end
    6097  : begin
              real_value= 30369;
              imag_value=12288;
            end
    6098  : begin
              real_value= 27240;
              imag_value=18200;
            end
    6099  : begin
              real_value= 22974;
              imag_value=23354;
            end
    6100  : begin
              real_value= 17752;
              imag_value=27534;
            end
    6101  : begin
              real_value= 11790;
              imag_value=30565;
            end
    6102  : begin
              real_value= 5336;
              imag_value=32323;
            end
    6103  : begin
              real_value= -1338;
              imag_value=32733;
            end
    6104  : begin
              real_value= -7959;
              imag_value=31779;
            end
    6105  : begin
              real_value= -14248;
              imag_value=29499;
            end
    6106  : begin
              real_value= -19943;
              imag_value=25990;
            end
    6107  : begin
              real_value= -24806;
              imag_value=21399;
            end
    6108  : begin
              real_value= -28636;
              imag_value=15914;
            end
    6109  : begin
              real_value= -31271;
              imag_value=9765;
            end
    6110  : begin
              real_value= -32603;
              imag_value=3210;
            end
    6111  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    6112  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    6113  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    6114  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    6115  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    6116  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    6117  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    6118  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    6119  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    6120  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    6121  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    6122  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    6123  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    6124  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    6125  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    6126  : begin
              real_value= 32743;
              imag_value=1070;
            end
    6127  : begin
              real_value= 31843;
              imag_value=7699;
            end
    6128  : begin
              real_value= 29615;
              imag_value=14006;
            end
    6129  : begin
              real_value= 26152;
              imag_value=19729;
            end
    6130  : begin
              real_value= 21600;
              imag_value=24630;
            end
    6131  : begin
              real_value= 16148;
              imag_value=28506;
            end
    6132  : begin
              real_value= 10021;
              imag_value=31191;
            end
    6133  : begin
              real_value= 3476;
              imag_value=32575;
            end
    6134  : begin
              real_value= -3210;
              imag_value=32603;
            end
    6135  : begin
              real_value= -9765;
              imag_value=31271;
            end
    6136  : begin
              real_value= -15914;
              imag_value=28636;
            end
    6137  : begin
              real_value= -21399;
              imag_value=24806;
            end
    6138  : begin
              real_value= -25990;
              imag_value=19943;
            end
    6139  : begin
              real_value= -29499;
              imag_value=14248;
            end
    6140  : begin
              real_value= -31779;
              imag_value=7959;
            end
    6141  : begin
              real_value= -32733;
              imag_value=1338;
            end
    6142  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    6143  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    6144  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    6145  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    6146  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    6147  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    6148  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    6149  : begin
              real_value= 802;
              imag_value=-32750;
            end
    6150  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    6151  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    6152  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    6153  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    6154  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    6155  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    6156  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    6157  : begin
              real_value= 32629;
              imag_value=2942;
            end
    6158  : begin
              real_value= 31351;
              imag_value=9508;
            end
    6159  : begin
              real_value= 28766;
              imag_value=15678;
            end
    6160  : begin
              real_value= 24981;
              imag_value=21194;
            end
    6161  : begin
              real_value= 20154;
              imag_value=25826;
            end
    6162  : begin
              real_value= 14489;
              imag_value=29382;
            end
    6163  : begin
              real_value= 8219;
              imag_value=31713;
            end
    6164  : begin
              real_value= 1606;
              imag_value=32721;
            end
    6165  : begin
              real_value= -5071;
              imag_value=32365;
            end
    6166  : begin
              real_value= -11539;
              imag_value=30661;
            end
    6167  : begin
              real_value= -17525;
              imag_value=27678;
            end
    6168  : begin
              real_value= -22782;
              imag_value=23541;
            end
    6169  : begin
              real_value= -27090;
              imag_value=18423;
            end
    6170  : begin
              real_value= -30267;
              imag_value=12537;
            end
    6171  : begin
              real_value= -32183;
              imag_value=6127;
            end
    6172  : begin
              real_value= -32757;
              imag_value=-535;
            end
    6173  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    6174  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    6175  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    6176  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    6177  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    6178  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    6179  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    6180  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    6181  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    6182  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    6183  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    6184  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    6185  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    6186  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    6187  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    6188  : begin
              real_value= 32407;
              imag_value=4806;
            end
    6189  : begin
              real_value= 30755;
              imag_value=11289;
            end
    6190  : begin
              real_value= 27820;
              imag_value=17299;
            end
    6191  : begin
              real_value= 23726;
              imag_value=22589;
            end
    6192  : begin
              real_value= 18644;
              imag_value=26938;
            end
    6193  : begin
              real_value= 12784;
              imag_value=30163;
            end
    6194  : begin
              real_value= 6390;
              imag_value=32131;
            end
    6195  : begin
              real_value= -267;
              imag_value=32759;
            end
    6196  : begin
              real_value= -6915;
              imag_value=32022;
            end
    6197  : begin
              real_value= -13274;
              imag_value=29950;
            end
    6198  : begin
              real_value= -19081;
              imag_value=26630;
            end
    6199  : begin
              real_value= -24092;
              imag_value=22199;
            end
    6200  : begin
              real_value= -28100;
              imag_value=16842;
            end
    6201  : begin
              real_value= -30935;
              imag_value=10783;
            end
    6202  : begin
              real_value= -32481;
              imag_value=4275;
            end
    6203  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    6204  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    6205  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    6206  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    6207  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    6208  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    6209  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    6210  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    6211  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    6212  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    6213  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    6214  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    6215  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    6216  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    6217  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    6218  : begin
              real_value= 32760;
              imag_value=0;
            end
    6219  : begin
              real_value= 32077;
              imag_value=6654;
            end
    6220  : begin
              real_value= 30057;
              imag_value=13030;
            end
    6221  : begin
              real_value= 26784;
              imag_value=18863;
            end
    6222  : begin
              real_value= 22395;
              imag_value=23911;
            end
    6223  : begin
              real_value= 17072;
              imag_value=27961;
            end
    6224  : begin
              real_value= 11036;
              imag_value=30846;
            end
    6225  : begin
              real_value= 4540;
              imag_value=32445;
            end
    6226  : begin
              real_value= -2142;
              imag_value=32691;
            end
    6227  : begin
              real_value= -8737;
              imag_value=31575;
            end
    6228  : begin
              real_value= -14968;
              imag_value=29142;
            end
    6229  : begin
              real_value= -20575;
              imag_value=25494;
            end
    6230  : begin
              real_value= -25324;
              imag_value=20783;
            end
    6231  : begin
              real_value= -29017;
              imag_value=15206;
            end
    6232  : begin
              real_value= -31501;
              imag_value=8995;
            end
    6233  : begin
              real_value= -32673;
              imag_value=2408;
            end
    6234  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    6235  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    6236  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    6237  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    6238  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    6239  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    6240  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    6241  : begin
              real_value= -267;
              imag_value=-32759;
            end
    6242  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    6243  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    6244  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    6245  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    6246  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    6247  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    6248  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    6249  : begin
              real_value= 32707;
              imag_value=1874;
            end
    6250  : begin
              real_value= 31645;
              imag_value=8477;
            end
    6251  : begin
              real_value= 29263;
              imag_value=14728;
            end
    6252  : begin
              real_value= 25661;
              imag_value=20365;
            end
    6253  : begin
              real_value= 20988;
              imag_value=25154;
            end
    6254  : begin
              real_value= 15442;
              imag_value=28892;
            end
    6255  : begin
              real_value= 9253;
              imag_value=31426;
            end
    6256  : begin
              real_value= 2676;
              imag_value=32651;
            end
    6257  : begin
              real_value= -4009;
              imag_value=32515;
            end
    6258  : begin
              real_value= -10529;
              imag_value=31023;
            end
    6259  : begin
              real_value= -16611;
              imag_value=28236;
            end
    6260  : begin
              real_value= -22001;
              imag_value=24274;
            end
    6261  : begin
              real_value= -26472;
              imag_value=19299;
            end
    6262  : begin
              real_value= -29841;
              imag_value=13520;
            end
    6263  : begin
              real_value= -31965;
              imag_value=7177;
            end
    6264  : begin
              real_value= -32757;
              imag_value=535;
            end
    6265  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    6266  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    6267  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    6268  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    6269  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    6270  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    6271  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    6272  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    6273  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    6274  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    6275  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    6276  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    6277  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    6278  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    6279  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    6280  : begin
              real_value= 32547;
              imag_value=3742;
            end
    6281  : begin
              real_value= 31107;
              imag_value=10275;
            end
    6282  : begin
              real_value= 28371;
              imag_value=16380;
            end
    6283  : begin
              real_value= 24453;
              imag_value=21801;
            end
    6284  : begin
              real_value= 19515;
              imag_value=26314;
            end
    6285  : begin
              real_value= 13764;
              imag_value=29729;
            end
    6286  : begin
              real_value= 7438;
              imag_value=31905;
            end
    6287  : begin
              real_value= 802;
              imag_value=32750;
            end
    6288  : begin
              real_value= -5864;
              imag_value=32231;
            end
    6289  : begin
              real_value= -12288;
              imag_value=30369;
            end
    6290  : begin
              real_value= -18200;
              imag_value=27240;
            end
    6291  : begin
              real_value= -23354;
              imag_value=22974;
            end
    6292  : begin
              real_value= -27534;
              imag_value=17752;
            end
    6293  : begin
              real_value= -30565;
              imag_value=11790;
            end
    6294  : begin
              real_value= -32323;
              imag_value=5336;
            end
    6295  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    6296  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    6297  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    6298  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    6299  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    6300  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    6301  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    6302  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    6303  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    6304  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    6305  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    6306  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    6307  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    6308  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    6309  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    6310  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    6311  : begin
              real_value= 32278;
              imag_value=5599;
            end
    6312  : begin
              real_value= 30468;
              imag_value=12039;
            end
    6313  : begin
              real_value= 27387;
              imag_value=17977;
            end
    6314  : begin
              real_value= 23165;
              imag_value=23165;
            end
    6315  : begin
              real_value= 17977;
              imag_value=27387;
            end
    6316  : begin
              real_value= 12039;
              imag_value=30468;
            end
    6317  : begin
              real_value= 5599;
              imag_value=32278;
            end
    6318  : begin
              real_value= -1070;
              imag_value=32743;
            end
    6319  : begin
              real_value= -7699;
              imag_value=31843;
            end
    6320  : begin
              real_value= -14006;
              imag_value=29615;
            end
    6321  : begin
              real_value= -19729;
              imag_value=26152;
            end
    6322  : begin
              real_value= -24630;
              imag_value=21600;
            end
    6323  : begin
              real_value= -28506;
              imag_value=16148;
            end
    6324  : begin
              real_value= -31191;
              imag_value=10021;
            end
    6325  : begin
              real_value= -32575;
              imag_value=3476;
            end
    6326  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    6327  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    6328  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    6329  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    6330  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    6331  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    6332  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    6333  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    6334  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    6335  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    6336  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    6337  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    6338  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    6339  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    6340  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    6341  : begin
              real_value= 32750;
              imag_value=802;
            end
    6342  : begin
              real_value= 31905;
              imag_value=7438;
            end
    6343  : begin
              real_value= 29729;
              imag_value=13764;
            end
    6344  : begin
              real_value= 26314;
              imag_value=19515;
            end
    6345  : begin
              real_value= 21801;
              imag_value=24453;
            end
    6346  : begin
              real_value= 16380;
              imag_value=28371;
            end
    6347  : begin
              real_value= 10275;
              imag_value=31107;
            end
    6348  : begin
              real_value= 3742;
              imag_value=32547;
            end
    6349  : begin
              real_value= -2942;
              imag_value=32629;
            end
    6350  : begin
              real_value= -9508;
              imag_value=31351;
            end
    6351  : begin
              real_value= -15678;
              imag_value=28766;
            end
    6352  : begin
              real_value= -21194;
              imag_value=24981;
            end
    6353  : begin
              real_value= -25826;
              imag_value=20154;
            end
    6354  : begin
              real_value= -29382;
              imag_value=14489;
            end
    6355  : begin
              real_value= -31713;
              imag_value=8219;
            end
    6356  : begin
              real_value= -32721;
              imag_value=1606;
            end
    6357  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    6358  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    6359  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    6360  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    6361  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    6362  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    6363  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    6364  : begin
              real_value= 535;
              imag_value=-32757;
            end
    6365  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    6366  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    6367  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    6368  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    6369  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    6370  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    6371  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    6372  : begin
              real_value= 32651;
              imag_value=2676;
            end
    6373  : begin
              real_value= 31426;
              imag_value=9253;
            end
    6374  : begin
              real_value= 28892;
              imag_value=15442;
            end
    6375  : begin
              real_value= 25154;
              imag_value=20988;
            end
    6376  : begin
              real_value= 20365;
              imag_value=25661;
            end
    6377  : begin
              real_value= 14728;
              imag_value=29263;
            end
    6378  : begin
              real_value= 8477;
              imag_value=31645;
            end
    6379  : begin
              real_value= 1874;
              imag_value=32707;
            end
    6380  : begin
              real_value= -4806;
              imag_value=32407;
            end
    6381  : begin
              real_value= -11289;
              imag_value=30755;
            end
    6382  : begin
              real_value= -17299;
              imag_value=27820;
            end
    6383  : begin
              real_value= -22589;
              imag_value=23726;
            end
    6384  : begin
              real_value= -26938;
              imag_value=18644;
            end
    6385  : begin
              real_value= -30163;
              imag_value=12784;
            end
    6386  : begin
              real_value= -32131;
              imag_value=6390;
            end
    6387  : begin
              real_value= -32759;
              imag_value=-267;
            end
    6388  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    6389  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    6390  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    6391  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    6392  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    6393  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    6394  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    6395  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    6396  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    6397  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    6398  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    6399  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    6400  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    6401  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    6402  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    6403  : begin
              real_value= 32445;
              imag_value=4540;
            end
    6404  : begin
              real_value= 30846;
              imag_value=11036;
            end
    6405  : begin
              real_value= 27961;
              imag_value=17072;
            end
    6406  : begin
              real_value= 23911;
              imag_value=22395;
            end
    6407  : begin
              real_value= 18863;
              imag_value=26784;
            end
    6408  : begin
              real_value= 13030;
              imag_value=30057;
            end
    6409  : begin
              real_value= 6654;
              imag_value=32077;
            end
    6410  : begin
              real_value= 0;
              imag_value=32760;
            end
    6411  : begin
              real_value= -6654;
              imag_value=32077;
            end
    6412  : begin
              real_value= -13030;
              imag_value=30057;
            end
    6413  : begin
              real_value= -18863;
              imag_value=26784;
            end
    6414  : begin
              real_value= -23911;
              imag_value=22395;
            end
    6415  : begin
              real_value= -27961;
              imag_value=17072;
            end
    6416  : begin
              real_value= -30846;
              imag_value=11036;
            end
    6417  : begin
              real_value= -32445;
              imag_value=4540;
            end
    6418  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    6419  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    6420  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    6421  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    6422  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    6423  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    6424  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    6425  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    6426  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    6427  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    6428  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    6429  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    6430  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    6431  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    6432  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    6433  : begin
              real_value= 32759;
              imag_value=-267;
            end
    6434  : begin
              real_value= 32131;
              imag_value=6390;
            end
    6435  : begin
              real_value= 30163;
              imag_value=12784;
            end
    6436  : begin
              real_value= 26938;
              imag_value=18644;
            end
    6437  : begin
              real_value= 22589;
              imag_value=23726;
            end
    6438  : begin
              real_value= 17299;
              imag_value=27820;
            end
    6439  : begin
              real_value= 11289;
              imag_value=30755;
            end
    6440  : begin
              real_value= 4806;
              imag_value=32407;
            end
    6441  : begin
              real_value= -1874;
              imag_value=32707;
            end
    6442  : begin
              real_value= -8477;
              imag_value=31645;
            end
    6443  : begin
              real_value= -14728;
              imag_value=29263;
            end
    6444  : begin
              real_value= -20365;
              imag_value=25661;
            end
    6445  : begin
              real_value= -25154;
              imag_value=20988;
            end
    6446  : begin
              real_value= -28892;
              imag_value=15442;
            end
    6447  : begin
              real_value= -31426;
              imag_value=9253;
            end
    6448  : begin
              real_value= -32651;
              imag_value=2676;
            end
    6449  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    6450  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    6451  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    6452  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    6453  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    6454  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    6455  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    6456  : begin
              real_value= -535;
              imag_value=-32757;
            end
    6457  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    6458  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    6459  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    6460  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    6461  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    6462  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    6463  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    6464  : begin
              real_value= 32721;
              imag_value=1606;
            end
    6465  : begin
              real_value= 31713;
              imag_value=8219;
            end
    6466  : begin
              real_value= 29382;
              imag_value=14489;
            end
    6467  : begin
              real_value= 25826;
              imag_value=20154;
            end
    6468  : begin
              real_value= 21194;
              imag_value=24981;
            end
    6469  : begin
              real_value= 15678;
              imag_value=28766;
            end
    6470  : begin
              real_value= 9508;
              imag_value=31351;
            end
    6471  : begin
              real_value= 2942;
              imag_value=32629;
            end
    6472  : begin
              real_value= -3742;
              imag_value=32547;
            end
    6473  : begin
              real_value= -10275;
              imag_value=31107;
            end
    6474  : begin
              real_value= -16380;
              imag_value=28371;
            end
    6475  : begin
              real_value= -21801;
              imag_value=24453;
            end
    6476  : begin
              real_value= -26314;
              imag_value=19515;
            end
    6477  : begin
              real_value= -29729;
              imag_value=13764;
            end
    6478  : begin
              real_value= -31905;
              imag_value=7438;
            end
    6479  : begin
              real_value= -32750;
              imag_value=802;
            end
    6480  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    6481  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    6482  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    6483  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    6484  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    6485  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    6486  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    6487  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    6488  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    6489  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    6490  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    6491  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    6492  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    6493  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    6494  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    6495  : begin
              real_value= 32575;
              imag_value=3476;
            end
    6496  : begin
              real_value= 31191;
              imag_value=10021;
            end
    6497  : begin
              real_value= 28506;
              imag_value=16148;
            end
    6498  : begin
              real_value= 24630;
              imag_value=21600;
            end
    6499  : begin
              real_value= 19729;
              imag_value=26152;
            end
    6500  : begin
              real_value= 14006;
              imag_value=29615;
            end
    6501  : begin
              real_value= 7699;
              imag_value=31843;
            end
    6502  : begin
              real_value= 1070;
              imag_value=32743;
            end
    6503  : begin
              real_value= -5599;
              imag_value=32278;
            end
    6504  : begin
              real_value= -12039;
              imag_value=30468;
            end
    6505  : begin
              real_value= -17977;
              imag_value=27387;
            end
    6506  : begin
              real_value= -23165;
              imag_value=23165;
            end
    6507  : begin
              real_value= -27387;
              imag_value=17977;
            end
    6508  : begin
              real_value= -30468;
              imag_value=12039;
            end
    6509  : begin
              real_value= -32278;
              imag_value=5599;
            end
    6510  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    6511  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    6512  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    6513  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    6514  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    6515  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    6516  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    6517  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    6518  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    6519  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    6520  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    6521  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    6522  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    6523  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    6524  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    6525  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    6526  : begin
              real_value= 32323;
              imag_value=5336;
            end
    6527  : begin
              real_value= 30565;
              imag_value=11790;
            end
    6528  : begin
              real_value= 27534;
              imag_value=17752;
            end
    6529  : begin
              real_value= 23354;
              imag_value=22974;
            end
    6530  : begin
              real_value= 18200;
              imag_value=27240;
            end
    6531  : begin
              real_value= 12288;
              imag_value=30369;
            end
    6532  : begin
              real_value= 5864;
              imag_value=32231;
            end
    6533  : begin
              real_value= -802;
              imag_value=32750;
            end
    6534  : begin
              real_value= -7438;
              imag_value=31905;
            end
    6535  : begin
              real_value= -13764;
              imag_value=29729;
            end
    6536  : begin
              real_value= -19515;
              imag_value=26314;
            end
    6537  : begin
              real_value= -24453;
              imag_value=21801;
            end
    6538  : begin
              real_value= -28371;
              imag_value=16380;
            end
    6539  : begin
              real_value= -31107;
              imag_value=10275;
            end
    6540  : begin
              real_value= -32547;
              imag_value=3742;
            end
    6541  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    6542  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    6543  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    6544  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    6545  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    6546  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    6547  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    6548  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    6549  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    6550  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    6551  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    6552  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    6553  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    6554  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    6555  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    6556  : begin
              real_value= 32757;
              imag_value=535;
            end
    6557  : begin
              real_value= 31965;
              imag_value=7177;
            end
    6558  : begin
              real_value= 29841;
              imag_value=13520;
            end
    6559  : begin
              real_value= 26472;
              imag_value=19299;
            end
    6560  : begin
              real_value= 22001;
              imag_value=24274;
            end
    6561  : begin
              real_value= 16611;
              imag_value=28236;
            end
    6562  : begin
              real_value= 10529;
              imag_value=31023;
            end
    6563  : begin
              real_value= 4009;
              imag_value=32515;
            end
    6564  : begin
              real_value= -2676;
              imag_value=32651;
            end
    6565  : begin
              real_value= -9253;
              imag_value=31426;
            end
    6566  : begin
              real_value= -15442;
              imag_value=28892;
            end
    6567  : begin
              real_value= -20988;
              imag_value=25154;
            end
    6568  : begin
              real_value= -25661;
              imag_value=20365;
            end
    6569  : begin
              real_value= -29263;
              imag_value=14728;
            end
    6570  : begin
              real_value= -31645;
              imag_value=8477;
            end
    6571  : begin
              real_value= -32707;
              imag_value=1874;
            end
    6572  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    6573  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    6574  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    6575  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    6576  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    6577  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    6578  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    6579  : begin
              real_value= 267;
              imag_value=-32759;
            end
    6580  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    6581  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    6582  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    6583  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    6584  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    6585  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    6586  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    6587  : begin
              real_value= 32673;
              imag_value=2408;
            end
    6588  : begin
              real_value= 31501;
              imag_value=8995;
            end
    6589  : begin
              real_value= 29017;
              imag_value=15206;
            end
    6590  : begin
              real_value= 25324;
              imag_value=20783;
            end
    6591  : begin
              real_value= 20575;
              imag_value=25494;
            end
    6592  : begin
              real_value= 14968;
              imag_value=29142;
            end
    6593  : begin
              real_value= 8737;
              imag_value=31575;
            end
    6594  : begin
              real_value= 2142;
              imag_value=32691;
            end
    6595  : begin
              real_value= -4540;
              imag_value=32445;
            end
    6596  : begin
              real_value= -11036;
              imag_value=30846;
            end
    6597  : begin
              real_value= -17072;
              imag_value=27961;
            end
    6598  : begin
              real_value= -22395;
              imag_value=23911;
            end
    6599  : begin
              real_value= -26784;
              imag_value=18863;
            end
    6600  : begin
              real_value= -30057;
              imag_value=13030;
            end
    6601  : begin
              real_value= -32077;
              imag_value=6654;
            end
    6602  : begin
              real_value= -32760;
              imag_value=0;
            end
    6603  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    6604  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    6605  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    6606  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    6607  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    6608  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    6609  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    6610  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    6611  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    6612  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    6613  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    6614  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    6615  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    6616  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    6617  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    6618  : begin
              real_value= 32481;
              imag_value=4275;
            end
    6619  : begin
              real_value= 30935;
              imag_value=10783;
            end
    6620  : begin
              real_value= 28100;
              imag_value=16842;
            end
    6621  : begin
              real_value= 24092;
              imag_value=22199;
            end
    6622  : begin
              real_value= 19081;
              imag_value=26630;
            end
    6623  : begin
              real_value= 13274;
              imag_value=29950;
            end
    6624  : begin
              real_value= 6915;
              imag_value=32022;
            end
    6625  : begin
              real_value= 267;
              imag_value=32759;
            end
    6626  : begin
              real_value= -6390;
              imag_value=32131;
            end
    6627  : begin
              real_value= -12784;
              imag_value=30163;
            end
    6628  : begin
              real_value= -18644;
              imag_value=26938;
            end
    6629  : begin
              real_value= -23726;
              imag_value=22589;
            end
    6630  : begin
              real_value= -27820;
              imag_value=17299;
            end
    6631  : begin
              real_value= -30755;
              imag_value=11289;
            end
    6632  : begin
              real_value= -32407;
              imag_value=4806;
            end
    6633  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    6634  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    6635  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    6636  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    6637  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    6638  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    6639  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    6640  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    6641  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    6642  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    6643  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    6644  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    6645  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    6646  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    6647  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    6648  : begin
              real_value= 32757;
              imag_value=-535;
            end
    6649  : begin
              real_value= 32183;
              imag_value=6127;
            end
    6650  : begin
              real_value= 30267;
              imag_value=12537;
            end
    6651  : begin
              real_value= 27090;
              imag_value=18423;
            end
    6652  : begin
              real_value= 22782;
              imag_value=23541;
            end
    6653  : begin
              real_value= 17525;
              imag_value=27678;
            end
    6654  : begin
              real_value= 11539;
              imag_value=30661;
            end
    6655  : begin
              real_value= 5071;
              imag_value=32365;
            end
    6656  : begin
              real_value= -1606;
              imag_value=32721;
            end
    6657  : begin
              real_value= -8219;
              imag_value=31713;
            end
    6658  : begin
              real_value= -14489;
              imag_value=29382;
            end
    6659  : begin
              real_value= -20154;
              imag_value=25826;
            end
    6660  : begin
              real_value= -24981;
              imag_value=21194;
            end
    6661  : begin
              real_value= -28766;
              imag_value=15678;
            end
    6662  : begin
              real_value= -31351;
              imag_value=9508;
            end
    6663  : begin
              real_value= -32629;
              imag_value=2942;
            end
    6664  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    6665  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    6666  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    6667  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    6668  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    6669  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    6670  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    6671  : begin
              real_value= -802;
              imag_value=-32750;
            end
    6672  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    6673  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    6674  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    6675  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    6676  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    6677  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    6678  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    6679  : begin
              real_value= 32733;
              imag_value=1338;
            end
    6680  : begin
              real_value= 31779;
              imag_value=7959;
            end
    6681  : begin
              real_value= 29499;
              imag_value=14248;
            end
    6682  : begin
              real_value= 25990;
              imag_value=19943;
            end
    6683  : begin
              real_value= 21399;
              imag_value=24806;
            end
    6684  : begin
              real_value= 15914;
              imag_value=28636;
            end
    6685  : begin
              real_value= 9765;
              imag_value=31271;
            end
    6686  : begin
              real_value= 3210;
              imag_value=32603;
            end
    6687  : begin
              real_value= -3476;
              imag_value=32575;
            end
    6688  : begin
              real_value= -10021;
              imag_value=31191;
            end
    6689  : begin
              real_value= -16148;
              imag_value=28506;
            end
    6690  : begin
              real_value= -21600;
              imag_value=24630;
            end
    6691  : begin
              real_value= -26152;
              imag_value=19729;
            end
    6692  : begin
              real_value= -29615;
              imag_value=14006;
            end
    6693  : begin
              real_value= -31843;
              imag_value=7699;
            end
    6694  : begin
              real_value= -32743;
              imag_value=1070;
            end
    6695  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    6696  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    6697  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    6698  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    6699  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    6700  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    6701  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    6702  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    6703  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    6704  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    6705  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    6706  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    6707  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    6708  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    6709  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    6710  : begin
              real_value= 32603;
              imag_value=3210;
            end
    6711  : begin
              real_value= 31271;
              imag_value=9765;
            end
    6712  : begin
              real_value= 28636;
              imag_value=15914;
            end
    6713  : begin
              real_value= 24806;
              imag_value=21399;
            end
    6714  : begin
              real_value= 19943;
              imag_value=25990;
            end
    6715  : begin
              real_value= 14248;
              imag_value=29499;
            end
    6716  : begin
              real_value= 7959;
              imag_value=31779;
            end
    6717  : begin
              real_value= 1338;
              imag_value=32733;
            end
    6718  : begin
              real_value= -5336;
              imag_value=32323;
            end
    6719  : begin
              real_value= -11790;
              imag_value=30565;
            end
    6720  : begin
              real_value= -17752;
              imag_value=27534;
            end
    6721  : begin
              real_value= -22974;
              imag_value=23354;
            end
    6722  : begin
              real_value= -27240;
              imag_value=18200;
            end
    6723  : begin
              real_value= -30369;
              imag_value=12288;
            end
    6724  : begin
              real_value= -32231;
              imag_value=5864;
            end
    6725  : begin
              real_value= -32750;
              imag_value=-802;
            end
    6726  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    6727  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    6728  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    6729  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    6730  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    6731  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    6732  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    6733  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    6734  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    6735  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    6736  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    6737  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    6738  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    6739  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    6740  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    6741  : begin
              real_value= 32365;
              imag_value=5071;
            end
    6742  : begin
              real_value= 30661;
              imag_value=11539;
            end
    6743  : begin
              real_value= 27678;
              imag_value=17525;
            end
    6744  : begin
              real_value= 23541;
              imag_value=22782;
            end
    6745  : begin
              real_value= 18423;
              imag_value=27090;
            end
    6746  : begin
              real_value= 12537;
              imag_value=30267;
            end
    6747  : begin
              real_value= 6127;
              imag_value=32183;
            end
    6748  : begin
              real_value= -535;
              imag_value=32757;
            end
    6749  : begin
              real_value= -7177;
              imag_value=31965;
            end
    6750  : begin
              real_value= -13520;
              imag_value=29841;
            end
    6751  : begin
              real_value= -19299;
              imag_value=26472;
            end
    6752  : begin
              real_value= -24274;
              imag_value=22001;
            end
    6753  : begin
              real_value= -28236;
              imag_value=16611;
            end
    6754  : begin
              real_value= -31023;
              imag_value=10529;
            end
    6755  : begin
              real_value= -32515;
              imag_value=4009;
            end
    6756  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    6757  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    6758  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    6759  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    6760  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    6761  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    6762  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    6763  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    6764  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    6765  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    6766  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    6767  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    6768  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    6769  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    6770  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    6771  : begin
              real_value= 32759;
              imag_value=267;
            end
    6772  : begin
              real_value= 32022;
              imag_value=6915;
            end
    6773  : begin
              real_value= 29950;
              imag_value=13274;
            end
    6774  : begin
              real_value= 26630;
              imag_value=19081;
            end
    6775  : begin
              real_value= 22199;
              imag_value=24092;
            end
    6776  : begin
              real_value= 16842;
              imag_value=28100;
            end
    6777  : begin
              real_value= 10783;
              imag_value=30935;
            end
    6778  : begin
              real_value= 4275;
              imag_value=32481;
            end
    6779  : begin
              real_value= -2408;
              imag_value=32673;
            end
    6780  : begin
              real_value= -8995;
              imag_value=31501;
            end
    6781  : begin
              real_value= -15206;
              imag_value=29017;
            end
    6782  : begin
              real_value= -20783;
              imag_value=25324;
            end
    6783  : begin
              real_value= -25494;
              imag_value=20575;
            end
    6784  : begin
              real_value= -29142;
              imag_value=14968;
            end
    6785  : begin
              real_value= -31575;
              imag_value=8737;
            end
    6786  : begin
              real_value= -32691;
              imag_value=2142;
            end
    6787  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    6788  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    6789  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    6790  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    6791  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    6792  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    6793  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    6794  : begin
              real_value= 0;
              imag_value=-32760;
            end
    6795  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    6796  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    6797  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    6798  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    6799  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    6800  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    6801  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    6802  : begin
              real_value= 32691;
              imag_value=2142;
            end
    6803  : begin
              real_value= 31575;
              imag_value=8737;
            end
    6804  : begin
              real_value= 29142;
              imag_value=14968;
            end
    6805  : begin
              real_value= 25494;
              imag_value=20575;
            end
    6806  : begin
              real_value= 20783;
              imag_value=25324;
            end
    6807  : begin
              real_value= 15206;
              imag_value=29017;
            end
    6808  : begin
              real_value= 8995;
              imag_value=31501;
            end
    6809  : begin
              real_value= 2408;
              imag_value=32673;
            end
    6810  : begin
              real_value= -4275;
              imag_value=32481;
            end
    6811  : begin
              real_value= -10783;
              imag_value=30935;
            end
    6812  : begin
              real_value= -16842;
              imag_value=28100;
            end
    6813  : begin
              real_value= -22199;
              imag_value=24092;
            end
    6814  : begin
              real_value= -26630;
              imag_value=19081;
            end
    6815  : begin
              real_value= -29950;
              imag_value=13274;
            end
    6816  : begin
              real_value= -32022;
              imag_value=6915;
            end
    6817  : begin
              real_value= -32759;
              imag_value=267;
            end
    6818  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    6819  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    6820  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    6821  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    6822  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    6823  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    6824  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    6825  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    6826  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    6827  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    6828  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    6829  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    6830  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    6831  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    6832  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    6833  : begin
              real_value= 32515;
              imag_value=4009;
            end
    6834  : begin
              real_value= 31023;
              imag_value=10529;
            end
    6835  : begin
              real_value= 28236;
              imag_value=16611;
            end
    6836  : begin
              real_value= 24274;
              imag_value=22001;
            end
    6837  : begin
              real_value= 19299;
              imag_value=26472;
            end
    6838  : begin
              real_value= 13520;
              imag_value=29841;
            end
    6839  : begin
              real_value= 7177;
              imag_value=31965;
            end
    6840  : begin
              real_value= 535;
              imag_value=32757;
            end
    6841  : begin
              real_value= -6127;
              imag_value=32183;
            end
    6842  : begin
              real_value= -12537;
              imag_value=30267;
            end
    6843  : begin
              real_value= -18423;
              imag_value=27090;
            end
    6844  : begin
              real_value= -23541;
              imag_value=22782;
            end
    6845  : begin
              real_value= -27678;
              imag_value=17525;
            end
    6846  : begin
              real_value= -30661;
              imag_value=11539;
            end
    6847  : begin
              real_value= -32365;
              imag_value=5071;
            end
    6848  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    6849  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    6850  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    6851  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    6852  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    6853  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    6854  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    6855  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    6856  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    6857  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    6858  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    6859  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    6860  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    6861  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    6862  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    6863  : begin
              real_value= 32750;
              imag_value=-802;
            end
    6864  : begin
              real_value= 32231;
              imag_value=5864;
            end
    6865  : begin
              real_value= 30369;
              imag_value=12288;
            end
    6866  : begin
              real_value= 27240;
              imag_value=18200;
            end
    6867  : begin
              real_value= 22974;
              imag_value=23354;
            end
    6868  : begin
              real_value= 17752;
              imag_value=27534;
            end
    6869  : begin
              real_value= 11790;
              imag_value=30565;
            end
    6870  : begin
              real_value= 5336;
              imag_value=32323;
            end
    6871  : begin
              real_value= -1338;
              imag_value=32733;
            end
    6872  : begin
              real_value= -7959;
              imag_value=31779;
            end
    6873  : begin
              real_value= -14248;
              imag_value=29499;
            end
    6874  : begin
              real_value= -19943;
              imag_value=25990;
            end
    6875  : begin
              real_value= -24806;
              imag_value=21399;
            end
    6876  : begin
              real_value= -28636;
              imag_value=15914;
            end
    6877  : begin
              real_value= -31271;
              imag_value=9765;
            end
    6878  : begin
              real_value= -32603;
              imag_value=3210;
            end
    6879  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    6880  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    6881  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    6882  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    6883  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    6884  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    6885  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    6886  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    6887  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    6888  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    6889  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    6890  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    6891  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    6892  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    6893  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    6894  : begin
              real_value= 32743;
              imag_value=1070;
            end
    6895  : begin
              real_value= 31843;
              imag_value=7699;
            end
    6896  : begin
              real_value= 29615;
              imag_value=14006;
            end
    6897  : begin
              real_value= 26152;
              imag_value=19729;
            end
    6898  : begin
              real_value= 21600;
              imag_value=24630;
            end
    6899  : begin
              real_value= 16148;
              imag_value=28506;
            end
    6900  : begin
              real_value= 10021;
              imag_value=31191;
            end
    6901  : begin
              real_value= 3476;
              imag_value=32575;
            end
    6902  : begin
              real_value= -3210;
              imag_value=32603;
            end
    6903  : begin
              real_value= -9765;
              imag_value=31271;
            end
    6904  : begin
              real_value= -15914;
              imag_value=28636;
            end
    6905  : begin
              real_value= -21399;
              imag_value=24806;
            end
    6906  : begin
              real_value= -25990;
              imag_value=19943;
            end
    6907  : begin
              real_value= -29499;
              imag_value=14248;
            end
    6908  : begin
              real_value= -31779;
              imag_value=7959;
            end
    6909  : begin
              real_value= -32733;
              imag_value=1338;
            end
    6910  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    6911  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    6912  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    6913  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    6914  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    6915  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    6916  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    6917  : begin
              real_value= 802;
              imag_value=-32750;
            end
    6918  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    6919  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    6920  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    6921  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    6922  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    6923  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    6924  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    6925  : begin
              real_value= 32629;
              imag_value=2942;
            end
    6926  : begin
              real_value= 31351;
              imag_value=9508;
            end
    6927  : begin
              real_value= 28766;
              imag_value=15678;
            end
    6928  : begin
              real_value= 24981;
              imag_value=21194;
            end
    6929  : begin
              real_value= 20154;
              imag_value=25826;
            end
    6930  : begin
              real_value= 14489;
              imag_value=29382;
            end
    6931  : begin
              real_value= 8219;
              imag_value=31713;
            end
    6932  : begin
              real_value= 1606;
              imag_value=32721;
            end
    6933  : begin
              real_value= -5071;
              imag_value=32365;
            end
    6934  : begin
              real_value= -11539;
              imag_value=30661;
            end
    6935  : begin
              real_value= -17525;
              imag_value=27678;
            end
    6936  : begin
              real_value= -22782;
              imag_value=23541;
            end
    6937  : begin
              real_value= -27090;
              imag_value=18423;
            end
    6938  : begin
              real_value= -30267;
              imag_value=12537;
            end
    6939  : begin
              real_value= -32183;
              imag_value=6127;
            end
    6940  : begin
              real_value= -32757;
              imag_value=-535;
            end
    6941  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    6942  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    6943  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    6944  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    6945  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    6946  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    6947  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    6948  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    6949  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    6950  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    6951  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    6952  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    6953  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    6954  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    6955  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    6956  : begin
              real_value= 32407;
              imag_value=4806;
            end
    6957  : begin
              real_value= 30755;
              imag_value=11289;
            end
    6958  : begin
              real_value= 27820;
              imag_value=17299;
            end
    6959  : begin
              real_value= 23726;
              imag_value=22589;
            end
    6960  : begin
              real_value= 18644;
              imag_value=26938;
            end
    6961  : begin
              real_value= 12784;
              imag_value=30163;
            end
    6962  : begin
              real_value= 6390;
              imag_value=32131;
            end
    6963  : begin
              real_value= -267;
              imag_value=32759;
            end
    6964  : begin
              real_value= -6915;
              imag_value=32022;
            end
    6965  : begin
              real_value= -13274;
              imag_value=29950;
            end
    6966  : begin
              real_value= -19081;
              imag_value=26630;
            end
    6967  : begin
              real_value= -24092;
              imag_value=22199;
            end
    6968  : begin
              real_value= -28100;
              imag_value=16842;
            end
    6969  : begin
              real_value= -30935;
              imag_value=10783;
            end
    6970  : begin
              real_value= -32481;
              imag_value=4275;
            end
    6971  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    6972  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    6973  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    6974  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    6975  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    6976  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    6977  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    6978  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    6979  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    6980  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    6981  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    6982  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    6983  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    6984  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    6985  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    6986  : begin
              real_value= 32760;
              imag_value=0;
            end
    6987  : begin
              real_value= 32077;
              imag_value=6654;
            end
    6988  : begin
              real_value= 30057;
              imag_value=13030;
            end
    6989  : begin
              real_value= 26784;
              imag_value=18863;
            end
    6990  : begin
              real_value= 22395;
              imag_value=23911;
            end
    6991  : begin
              real_value= 17072;
              imag_value=27961;
            end
    6992  : begin
              real_value= 11036;
              imag_value=30846;
            end
    6993  : begin
              real_value= 4540;
              imag_value=32445;
            end
    6994  : begin
              real_value= -2142;
              imag_value=32691;
            end
    6995  : begin
              real_value= -8737;
              imag_value=31575;
            end
    6996  : begin
              real_value= -14968;
              imag_value=29142;
            end
    6997  : begin
              real_value= -20575;
              imag_value=25494;
            end
    6998  : begin
              real_value= -25324;
              imag_value=20783;
            end
    6999  : begin
              real_value= -29017;
              imag_value=15206;
            end
    7000  : begin
              real_value= -31501;
              imag_value=8995;
            end
    7001  : begin
              real_value= -32673;
              imag_value=2408;
            end
    7002  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    7003  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    7004  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    7005  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    7006  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    7007  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    7008  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    7009  : begin
              real_value= -267;
              imag_value=-32759;
            end
    7010  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    7011  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    7012  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    7013  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    7014  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    7015  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    7016  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    7017  : begin
              real_value= 32707;
              imag_value=1874;
            end
    7018  : begin
              real_value= 31645;
              imag_value=8477;
            end
    7019  : begin
              real_value= 29263;
              imag_value=14728;
            end
    7020  : begin
              real_value= 25661;
              imag_value=20365;
            end
    7021  : begin
              real_value= 20988;
              imag_value=25154;
            end
    7022  : begin
              real_value= 15442;
              imag_value=28892;
            end
    7023  : begin
              real_value= 9253;
              imag_value=31426;
            end
    7024  : begin
              real_value= 2676;
              imag_value=32651;
            end
    7025  : begin
              real_value= -4009;
              imag_value=32515;
            end
    7026  : begin
              real_value= -10529;
              imag_value=31023;
            end
    7027  : begin
              real_value= -16611;
              imag_value=28236;
            end
    7028  : begin
              real_value= -22001;
              imag_value=24274;
            end
    7029  : begin
              real_value= -26472;
              imag_value=19299;
            end
    7030  : begin
              real_value= -29841;
              imag_value=13520;
            end
    7031  : begin
              real_value= -31965;
              imag_value=7177;
            end
    7032  : begin
              real_value= -32757;
              imag_value=535;
            end
    7033  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    7034  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    7035  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    7036  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    7037  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    7038  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    7039  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    7040  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    7041  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    7042  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    7043  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    7044  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    7045  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    7046  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    7047  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    7048  : begin
              real_value= 32547;
              imag_value=3742;
            end
    7049  : begin
              real_value= 31107;
              imag_value=10275;
            end
    7050  : begin
              real_value= 28371;
              imag_value=16380;
            end
    7051  : begin
              real_value= 24453;
              imag_value=21801;
            end
    7052  : begin
              real_value= 19515;
              imag_value=26314;
            end
    7053  : begin
              real_value= 13764;
              imag_value=29729;
            end
    7054  : begin
              real_value= 7438;
              imag_value=31905;
            end
    7055  : begin
              real_value= 802;
              imag_value=32750;
            end
    7056  : begin
              real_value= -5864;
              imag_value=32231;
            end
    7057  : begin
              real_value= -12288;
              imag_value=30369;
            end
    7058  : begin
              real_value= -18200;
              imag_value=27240;
            end
    7059  : begin
              real_value= -23354;
              imag_value=22974;
            end
    7060  : begin
              real_value= -27534;
              imag_value=17752;
            end
    7061  : begin
              real_value= -30565;
              imag_value=11790;
            end
    7062  : begin
              real_value= -32323;
              imag_value=5336;
            end
    7063  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    7064  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    7065  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    7066  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    7067  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    7068  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    7069  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    7070  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    7071  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    7072  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    7073  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    7074  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    7075  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    7076  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    7077  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    7078  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    7079  : begin
              real_value= 32278;
              imag_value=5599;
            end
    7080  : begin
              real_value= 30468;
              imag_value=12039;
            end
    7081  : begin
              real_value= 27387;
              imag_value=17977;
            end
    7082  : begin
              real_value= 23165;
              imag_value=23165;
            end
    7083  : begin
              real_value= 17977;
              imag_value=27387;
            end
    7084  : begin
              real_value= 12039;
              imag_value=30468;
            end
    7085  : begin
              real_value= 5599;
              imag_value=32278;
            end
    7086  : begin
              real_value= -1070;
              imag_value=32743;
            end
    7087  : begin
              real_value= -7699;
              imag_value=31843;
            end
    7088  : begin
              real_value= -14006;
              imag_value=29615;
            end
    7089  : begin
              real_value= -19729;
              imag_value=26152;
            end
    7090  : begin
              real_value= -24630;
              imag_value=21600;
            end
    7091  : begin
              real_value= -28506;
              imag_value=16148;
            end
    7092  : begin
              real_value= -31191;
              imag_value=10021;
            end
    7093  : begin
              real_value= -32575;
              imag_value=3476;
            end
    7094  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    7095  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    7096  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    7097  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    7098  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    7099  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    7100  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    7101  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    7102  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    7103  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    7104  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    7105  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    7106  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    7107  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    7108  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    7109  : begin
              real_value= 32750;
              imag_value=802;
            end
    7110  : begin
              real_value= 31905;
              imag_value=7438;
            end
    7111  : begin
              real_value= 29729;
              imag_value=13764;
            end
    7112  : begin
              real_value= 26314;
              imag_value=19515;
            end
    7113  : begin
              real_value= 21801;
              imag_value=24453;
            end
    7114  : begin
              real_value= 16380;
              imag_value=28371;
            end
    7115  : begin
              real_value= 10275;
              imag_value=31107;
            end
    7116  : begin
              real_value= 3742;
              imag_value=32547;
            end
    7117  : begin
              real_value= -2942;
              imag_value=32629;
            end
    7118  : begin
              real_value= -9508;
              imag_value=31351;
            end
    7119  : begin
              real_value= -15678;
              imag_value=28766;
            end
    7120  : begin
              real_value= -21194;
              imag_value=24981;
            end
    7121  : begin
              real_value= -25826;
              imag_value=20154;
            end
    7122  : begin
              real_value= -29382;
              imag_value=14489;
            end
    7123  : begin
              real_value= -31713;
              imag_value=8219;
            end
    7124  : begin
              real_value= -32721;
              imag_value=1606;
            end
    7125  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    7126  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    7127  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    7128  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    7129  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    7130  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    7131  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    7132  : begin
              real_value= 535;
              imag_value=-32757;
            end
    7133  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    7134  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    7135  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    7136  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    7137  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    7138  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    7139  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    7140  : begin
              real_value= 32651;
              imag_value=2676;
            end
    7141  : begin
              real_value= 31426;
              imag_value=9253;
            end
    7142  : begin
              real_value= 28892;
              imag_value=15442;
            end
    7143  : begin
              real_value= 25154;
              imag_value=20988;
            end
    7144  : begin
              real_value= 20365;
              imag_value=25661;
            end
    7145  : begin
              real_value= 14728;
              imag_value=29263;
            end
    7146  : begin
              real_value= 8477;
              imag_value=31645;
            end
    7147  : begin
              real_value= 1874;
              imag_value=32707;
            end
    7148  : begin
              real_value= -4806;
              imag_value=32407;
            end
    7149  : begin
              real_value= -11289;
              imag_value=30755;
            end
    7150  : begin
              real_value= -17299;
              imag_value=27820;
            end
    7151  : begin
              real_value= -22589;
              imag_value=23726;
            end
    7152  : begin
              real_value= -26938;
              imag_value=18644;
            end
    7153  : begin
              real_value= -30163;
              imag_value=12784;
            end
    7154  : begin
              real_value= -32131;
              imag_value=6390;
            end
    7155  : begin
              real_value= -32759;
              imag_value=-267;
            end
    7156  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    7157  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    7158  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    7159  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    7160  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    7161  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    7162  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    7163  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    7164  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    7165  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    7166  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    7167  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    7168  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    7169  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    7170  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    7171  : begin
              real_value= 32445;
              imag_value=4540;
            end
    7172  : begin
              real_value= 30846;
              imag_value=11036;
            end
    7173  : begin
              real_value= 27961;
              imag_value=17072;
            end
    7174  : begin
              real_value= 23911;
              imag_value=22395;
            end
    7175  : begin
              real_value= 18863;
              imag_value=26784;
            end
    7176  : begin
              real_value= 13030;
              imag_value=30057;
            end
    7177  : begin
              real_value= 6654;
              imag_value=32077;
            end
    7178  : begin
              real_value= 0;
              imag_value=32760;
            end
    7179  : begin
              real_value= -6654;
              imag_value=32077;
            end
    7180  : begin
              real_value= -13030;
              imag_value=30057;
            end
    7181  : begin
              real_value= -18863;
              imag_value=26784;
            end
    7182  : begin
              real_value= -23911;
              imag_value=22395;
            end
    7183  : begin
              real_value= -27961;
              imag_value=17072;
            end
    7184  : begin
              real_value= -30846;
              imag_value=11036;
            end
    7185  : begin
              real_value= -32445;
              imag_value=4540;
            end
    7186  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    7187  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    7188  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    7189  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    7190  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    7191  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    7192  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    7193  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    7194  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    7195  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    7196  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    7197  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    7198  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    7199  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    7200  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    7201  : begin
              real_value= 32759;
              imag_value=-267;
            end
    7202  : begin
              real_value= 32131;
              imag_value=6390;
            end
    7203  : begin
              real_value= 30163;
              imag_value=12784;
            end
    7204  : begin
              real_value= 26938;
              imag_value=18644;
            end
    7205  : begin
              real_value= 22589;
              imag_value=23726;
            end
    7206  : begin
              real_value= 17299;
              imag_value=27820;
            end
    7207  : begin
              real_value= 11289;
              imag_value=30755;
            end
    7208  : begin
              real_value= 4806;
              imag_value=32407;
            end
    7209  : begin
              real_value= -1874;
              imag_value=32707;
            end
    7210  : begin
              real_value= -8477;
              imag_value=31645;
            end
    7211  : begin
              real_value= -14728;
              imag_value=29263;
            end
    7212  : begin
              real_value= -20365;
              imag_value=25661;
            end
    7213  : begin
              real_value= -25154;
              imag_value=20988;
            end
    7214  : begin
              real_value= -28892;
              imag_value=15442;
            end
    7215  : begin
              real_value= -31426;
              imag_value=9253;
            end
    7216  : begin
              real_value= -32651;
              imag_value=2676;
            end
    7217  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    7218  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    7219  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    7220  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    7221  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    7222  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    7223  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    7224  : begin
              real_value= -535;
              imag_value=-32757;
            end
    7225  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    7226  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    7227  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    7228  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    7229  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    7230  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    7231  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    7232  : begin
              real_value= 32721;
              imag_value=1606;
            end
    7233  : begin
              real_value= 31713;
              imag_value=8219;
            end
    7234  : begin
              real_value= 29382;
              imag_value=14489;
            end
    7235  : begin
              real_value= 25826;
              imag_value=20154;
            end
    7236  : begin
              real_value= 21194;
              imag_value=24981;
            end
    7237  : begin
              real_value= 15678;
              imag_value=28766;
            end
    7238  : begin
              real_value= 9508;
              imag_value=31351;
            end
    7239  : begin
              real_value= 2942;
              imag_value=32629;
            end
    7240  : begin
              real_value= -3742;
              imag_value=32547;
            end
    7241  : begin
              real_value= -10275;
              imag_value=31107;
            end
    7242  : begin
              real_value= -16380;
              imag_value=28371;
            end
    7243  : begin
              real_value= -21801;
              imag_value=24453;
            end
    7244  : begin
              real_value= -26314;
              imag_value=19515;
            end
    7245  : begin
              real_value= -29729;
              imag_value=13764;
            end
    7246  : begin
              real_value= -31905;
              imag_value=7438;
            end
    7247  : begin
              real_value= -32750;
              imag_value=802;
            end
    7248  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    7249  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    7250  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    7251  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    7252  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    7253  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    7254  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    7255  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    7256  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    7257  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    7258  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    7259  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    7260  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    7261  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    7262  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    7263  : begin
              real_value= 32575;
              imag_value=3476;
            end
    7264  : begin
              real_value= 31191;
              imag_value=10021;
            end
    7265  : begin
              real_value= 28506;
              imag_value=16148;
            end
    7266  : begin
              real_value= 24630;
              imag_value=21600;
            end
    7267  : begin
              real_value= 19729;
              imag_value=26152;
            end
    7268  : begin
              real_value= 14006;
              imag_value=29615;
            end
    7269  : begin
              real_value= 7699;
              imag_value=31843;
            end
    7270  : begin
              real_value= 1070;
              imag_value=32743;
            end
    7271  : begin
              real_value= -5599;
              imag_value=32278;
            end
    7272  : begin
              real_value= -12039;
              imag_value=30468;
            end
    7273  : begin
              real_value= -17977;
              imag_value=27387;
            end
    7274  : begin
              real_value= -23165;
              imag_value=23165;
            end
    7275  : begin
              real_value= -27387;
              imag_value=17977;
            end
    7276  : begin
              real_value= -30468;
              imag_value=12039;
            end
    7277  : begin
              real_value= -32278;
              imag_value=5599;
            end
    7278  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    7279  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    7280  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    7281  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    7282  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    7283  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    7284  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    7285  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    7286  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    7287  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    7288  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    7289  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    7290  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    7291  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    7292  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    7293  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    7294  : begin
              real_value= 32323;
              imag_value=5336;
            end
    7295  : begin
              real_value= 30565;
              imag_value=11790;
            end
    7296  : begin
              real_value= 27534;
              imag_value=17752;
            end
    7297  : begin
              real_value= 23354;
              imag_value=22974;
            end
    7298  : begin
              real_value= 18200;
              imag_value=27240;
            end
    7299  : begin
              real_value= 12288;
              imag_value=30369;
            end
    7300  : begin
              real_value= 5864;
              imag_value=32231;
            end
    7301  : begin
              real_value= -802;
              imag_value=32750;
            end
    7302  : begin
              real_value= -7438;
              imag_value=31905;
            end
    7303  : begin
              real_value= -13764;
              imag_value=29729;
            end
    7304  : begin
              real_value= -19515;
              imag_value=26314;
            end
    7305  : begin
              real_value= -24453;
              imag_value=21801;
            end
    7306  : begin
              real_value= -28371;
              imag_value=16380;
            end
    7307  : begin
              real_value= -31107;
              imag_value=10275;
            end
    7308  : begin
              real_value= -32547;
              imag_value=3742;
            end
    7309  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    7310  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    7311  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    7312  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    7313  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    7314  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    7315  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    7316  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    7317  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    7318  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    7319  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    7320  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    7321  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    7322  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    7323  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    7324  : begin
              real_value= 32757;
              imag_value=535;
            end
    7325  : begin
              real_value= 31965;
              imag_value=7177;
            end
    7326  : begin
              real_value= 29841;
              imag_value=13520;
            end
    7327  : begin
              real_value= 26472;
              imag_value=19299;
            end
    7328  : begin
              real_value= 22001;
              imag_value=24274;
            end
    7329  : begin
              real_value= 16611;
              imag_value=28236;
            end
    7330  : begin
              real_value= 10529;
              imag_value=31023;
            end
    7331  : begin
              real_value= 4009;
              imag_value=32515;
            end
    7332  : begin
              real_value= -2676;
              imag_value=32651;
            end
    7333  : begin
              real_value= -9253;
              imag_value=31426;
            end
    7334  : begin
              real_value= -15442;
              imag_value=28892;
            end
    7335  : begin
              real_value= -20988;
              imag_value=25154;
            end
    7336  : begin
              real_value= -25661;
              imag_value=20365;
            end
    7337  : begin
              real_value= -29263;
              imag_value=14728;
            end
    7338  : begin
              real_value= -31645;
              imag_value=8477;
            end
    7339  : begin
              real_value= -32707;
              imag_value=1874;
            end
    7340  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    7341  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    7342  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    7343  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    7344  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    7345  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    7346  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    7347  : begin
              real_value= 267;
              imag_value=-32759;
            end
    7348  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    7349  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    7350  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    7351  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    7352  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    7353  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    7354  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    7355  : begin
              real_value= 32673;
              imag_value=2408;
            end
    7356  : begin
              real_value= 31501;
              imag_value=8995;
            end
    7357  : begin
              real_value= 29017;
              imag_value=15206;
            end
    7358  : begin
              real_value= 25324;
              imag_value=20783;
            end
    7359  : begin
              real_value= 20575;
              imag_value=25494;
            end
    7360  : begin
              real_value= 14968;
              imag_value=29142;
            end
    7361  : begin
              real_value= 8737;
              imag_value=31575;
            end
    7362  : begin
              real_value= 2142;
              imag_value=32691;
            end
    7363  : begin
              real_value= -4540;
              imag_value=32445;
            end
    7364  : begin
              real_value= -11036;
              imag_value=30846;
            end
    7365  : begin
              real_value= -17072;
              imag_value=27961;
            end
    7366  : begin
              real_value= -22395;
              imag_value=23911;
            end
    7367  : begin
              real_value= -26784;
              imag_value=18863;
            end
    7368  : begin
              real_value= -30057;
              imag_value=13030;
            end
    7369  : begin
              real_value= -32077;
              imag_value=6654;
            end
    7370  : begin
              real_value= -32760;
              imag_value=0;
            end
    7371  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    7372  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    7373  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    7374  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    7375  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    7376  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    7377  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    7378  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    7379  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    7380  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    7381  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    7382  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    7383  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    7384  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    7385  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    7386  : begin
              real_value= 32481;
              imag_value=4275;
            end
    7387  : begin
              real_value= 30935;
              imag_value=10783;
            end
    7388  : begin
              real_value= 28100;
              imag_value=16842;
            end
    7389  : begin
              real_value= 24092;
              imag_value=22199;
            end
    7390  : begin
              real_value= 19081;
              imag_value=26630;
            end
    7391  : begin
              real_value= 13274;
              imag_value=29950;
            end
    7392  : begin
              real_value= 6915;
              imag_value=32022;
            end
    7393  : begin
              real_value= 267;
              imag_value=32759;
            end
    7394  : begin
              real_value= -6390;
              imag_value=32131;
            end
    7395  : begin
              real_value= -12784;
              imag_value=30163;
            end
    7396  : begin
              real_value= -18644;
              imag_value=26938;
            end
    7397  : begin
              real_value= -23726;
              imag_value=22589;
            end
    7398  : begin
              real_value= -27820;
              imag_value=17299;
            end
    7399  : begin
              real_value= -30755;
              imag_value=11289;
            end
    7400  : begin
              real_value= -32407;
              imag_value=4806;
            end
    7401  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    7402  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    7403  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    7404  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    7405  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    7406  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    7407  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    7408  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    7409  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    7410  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    7411  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    7412  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    7413  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    7414  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    7415  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    7416  : begin
              real_value= 32757;
              imag_value=-535;
            end
    7417  : begin
              real_value= 32183;
              imag_value=6127;
            end
    7418  : begin
              real_value= 30267;
              imag_value=12537;
            end
    7419  : begin
              real_value= 27090;
              imag_value=18423;
            end
    7420  : begin
              real_value= 22782;
              imag_value=23541;
            end
    7421  : begin
              real_value= 17525;
              imag_value=27678;
            end
    7422  : begin
              real_value= 11539;
              imag_value=30661;
            end
    7423  : begin
              real_value= 5071;
              imag_value=32365;
            end
    7424  : begin
              real_value= -1606;
              imag_value=32721;
            end
    7425  : begin
              real_value= -8219;
              imag_value=31713;
            end
    7426  : begin
              real_value= -14489;
              imag_value=29382;
            end
    7427  : begin
              real_value= -20154;
              imag_value=25826;
            end
    7428  : begin
              real_value= -24981;
              imag_value=21194;
            end
    7429  : begin
              real_value= -28766;
              imag_value=15678;
            end
    7430  : begin
              real_value= -31351;
              imag_value=9508;
            end
    7431  : begin
              real_value= -32629;
              imag_value=2942;
            end
    7432  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    7433  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    7434  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    7435  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    7436  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    7437  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    7438  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    7439  : begin
              real_value= -802;
              imag_value=-32750;
            end
    7440  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    7441  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    7442  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    7443  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    7444  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    7445  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    7446  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    7447  : begin
              real_value= 32733;
              imag_value=1338;
            end
    7448  : begin
              real_value= 31779;
              imag_value=7959;
            end
    7449  : begin
              real_value= 29499;
              imag_value=14248;
            end
    7450  : begin
              real_value= 25990;
              imag_value=19943;
            end
    7451  : begin
              real_value= 21399;
              imag_value=24806;
            end
    7452  : begin
              real_value= 15914;
              imag_value=28636;
            end
    7453  : begin
              real_value= 9765;
              imag_value=31271;
            end
    7454  : begin
              real_value= 3210;
              imag_value=32603;
            end
    7455  : begin
              real_value= -3476;
              imag_value=32575;
            end
    7456  : begin
              real_value= -10021;
              imag_value=31191;
            end
    7457  : begin
              real_value= -16148;
              imag_value=28506;
            end
    7458  : begin
              real_value= -21600;
              imag_value=24630;
            end
    7459  : begin
              real_value= -26152;
              imag_value=19729;
            end
    7460  : begin
              real_value= -29615;
              imag_value=14006;
            end
    7461  : begin
              real_value= -31843;
              imag_value=7699;
            end
    7462  : begin
              real_value= -32743;
              imag_value=1070;
            end
    7463  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    7464  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    7465  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    7466  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    7467  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    7468  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    7469  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    7470  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    7471  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    7472  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    7473  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    7474  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    7475  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    7476  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    7477  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    7478  : begin
              real_value= 32603;
              imag_value=3210;
            end
    7479  : begin
              real_value= 31271;
              imag_value=9765;
            end
    7480  : begin
              real_value= 28636;
              imag_value=15914;
            end
    7481  : begin
              real_value= 24806;
              imag_value=21399;
            end
    7482  : begin
              real_value= 19943;
              imag_value=25990;
            end
    7483  : begin
              real_value= 14248;
              imag_value=29499;
            end
    7484  : begin
              real_value= 7959;
              imag_value=31779;
            end
    7485  : begin
              real_value= 1338;
              imag_value=32733;
            end
    7486  : begin
              real_value= -5336;
              imag_value=32323;
            end
    7487  : begin
              real_value= -11790;
              imag_value=30565;
            end
    7488  : begin
              real_value= -17752;
              imag_value=27534;
            end
    7489  : begin
              real_value= -22974;
              imag_value=23354;
            end
    7490  : begin
              real_value= -27240;
              imag_value=18200;
            end
    7491  : begin
              real_value= -30369;
              imag_value=12288;
            end
    7492  : begin
              real_value= -32231;
              imag_value=5864;
            end
    7493  : begin
              real_value= -32750;
              imag_value=-802;
            end
    7494  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    7495  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    7496  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    7497  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    7498  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    7499  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    7500  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    7501  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    7502  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    7503  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    7504  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    7505  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    7506  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    7507  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    7508  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    7509  : begin
              real_value= 32365;
              imag_value=5071;
            end
    7510  : begin
              real_value= 30661;
              imag_value=11539;
            end
    7511  : begin
              real_value= 27678;
              imag_value=17525;
            end
    7512  : begin
              real_value= 23541;
              imag_value=22782;
            end
    7513  : begin
              real_value= 18423;
              imag_value=27090;
            end
    7514  : begin
              real_value= 12537;
              imag_value=30267;
            end
    7515  : begin
              real_value= 6127;
              imag_value=32183;
            end
    7516  : begin
              real_value= -535;
              imag_value=32757;
            end
    7517  : begin
              real_value= -7177;
              imag_value=31965;
            end
    7518  : begin
              real_value= -13520;
              imag_value=29841;
            end
    7519  : begin
              real_value= -19299;
              imag_value=26472;
            end
    7520  : begin
              real_value= -24274;
              imag_value=22001;
            end
    7521  : begin
              real_value= -28236;
              imag_value=16611;
            end
    7522  : begin
              real_value= -31023;
              imag_value=10529;
            end
    7523  : begin
              real_value= -32515;
              imag_value=4009;
            end
    7524  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    7525  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    7526  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    7527  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    7528  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    7529  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    7530  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    7531  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    7532  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    7533  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    7534  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    7535  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    7536  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    7537  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    7538  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    7539  : begin
              real_value= 32759;
              imag_value=267;
            end
    7540  : begin
              real_value= 32022;
              imag_value=6915;
            end
    7541  : begin
              real_value= 29950;
              imag_value=13274;
            end
    7542  : begin
              real_value= 26630;
              imag_value=19081;
            end
    7543  : begin
              real_value= 22199;
              imag_value=24092;
            end
    7544  : begin
              real_value= 16842;
              imag_value=28100;
            end
    7545  : begin
              real_value= 10783;
              imag_value=30935;
            end
    7546  : begin
              real_value= 4275;
              imag_value=32481;
            end
    7547  : begin
              real_value= -2408;
              imag_value=32673;
            end
    7548  : begin
              real_value= -8995;
              imag_value=31501;
            end
    7549  : begin
              real_value= -15206;
              imag_value=29017;
            end
    7550  : begin
              real_value= -20783;
              imag_value=25324;
            end
    7551  : begin
              real_value= -25494;
              imag_value=20575;
            end
    7552  : begin
              real_value= -29142;
              imag_value=14968;
            end
    7553  : begin
              real_value= -31575;
              imag_value=8737;
            end
    7554  : begin
              real_value= -32691;
              imag_value=2142;
            end
    7555  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    7556  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    7557  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    7558  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    7559  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    7560  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    7561  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    7562  : begin
              real_value= 0;
              imag_value=-32760;
            end
    7563  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    7564  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    7565  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    7566  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    7567  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    7568  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    7569  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    7570  : begin
              real_value= 32691;
              imag_value=2142;
            end
    7571  : begin
              real_value= 31575;
              imag_value=8737;
            end
    7572  : begin
              real_value= 29142;
              imag_value=14968;
            end
    7573  : begin
              real_value= 25494;
              imag_value=20575;
            end
    7574  : begin
              real_value= 20783;
              imag_value=25324;
            end
    7575  : begin
              real_value= 15206;
              imag_value=29017;
            end
    7576  : begin
              real_value= 8995;
              imag_value=31501;
            end
    7577  : begin
              real_value= 2408;
              imag_value=32673;
            end
    7578  : begin
              real_value= -4275;
              imag_value=32481;
            end
    7579  : begin
              real_value= -10783;
              imag_value=30935;
            end
    7580  : begin
              real_value= -16842;
              imag_value=28100;
            end
    7581  : begin
              real_value= -22199;
              imag_value=24092;
            end
    7582  : begin
              real_value= -26630;
              imag_value=19081;
            end
    7583  : begin
              real_value= -29950;
              imag_value=13274;
            end
    7584  : begin
              real_value= -32022;
              imag_value=6915;
            end
    7585  : begin
              real_value= -32759;
              imag_value=267;
            end
    7586  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    7587  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    7588  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    7589  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    7590  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    7591  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    7592  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    7593  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    7594  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    7595  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    7596  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    7597  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    7598  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    7599  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    7600  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    7601  : begin
              real_value= 32515;
              imag_value=4009;
            end
    7602  : begin
              real_value= 31023;
              imag_value=10529;
            end
    7603  : begin
              real_value= 28236;
              imag_value=16611;
            end
    7604  : begin
              real_value= 24274;
              imag_value=22001;
            end
    7605  : begin
              real_value= 19299;
              imag_value=26472;
            end
    7606  : begin
              real_value= 13520;
              imag_value=29841;
            end
    7607  : begin
              real_value= 7177;
              imag_value=31965;
            end
    7608  : begin
              real_value= 535;
              imag_value=32757;
            end
    7609  : begin
              real_value= -6127;
              imag_value=32183;
            end
    7610  : begin
              real_value= -12537;
              imag_value=30267;
            end
    7611  : begin
              real_value= -18423;
              imag_value=27090;
            end
    7612  : begin
              real_value= -23541;
              imag_value=22782;
            end
    7613  : begin
              real_value= -27678;
              imag_value=17525;
            end
    7614  : begin
              real_value= -30661;
              imag_value=11539;
            end
    7615  : begin
              real_value= -32365;
              imag_value=5071;
            end
    7616  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    7617  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    7618  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    7619  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    7620  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    7621  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    7622  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    7623  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    7624  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    7625  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    7626  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    7627  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    7628  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    7629  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    7630  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    7631  : begin
              real_value= 32750;
              imag_value=-802;
            end
    7632  : begin
              real_value= 32231;
              imag_value=5864;
            end
    7633  : begin
              real_value= 30369;
              imag_value=12288;
            end
    7634  : begin
              real_value= 27240;
              imag_value=18200;
            end
    7635  : begin
              real_value= 22974;
              imag_value=23354;
            end
    7636  : begin
              real_value= 17752;
              imag_value=27534;
            end
    7637  : begin
              real_value= 11790;
              imag_value=30565;
            end
    7638  : begin
              real_value= 5336;
              imag_value=32323;
            end
    7639  : begin
              real_value= -1338;
              imag_value=32733;
            end
    7640  : begin
              real_value= -7959;
              imag_value=31779;
            end
    7641  : begin
              real_value= -14248;
              imag_value=29499;
            end
    7642  : begin
              real_value= -19943;
              imag_value=25990;
            end
    7643  : begin
              real_value= -24806;
              imag_value=21399;
            end
    7644  : begin
              real_value= -28636;
              imag_value=15914;
            end
    7645  : begin
              real_value= -31271;
              imag_value=9765;
            end
    7646  : begin
              real_value= -32603;
              imag_value=3210;
            end
    7647  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    7648  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    7649  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    7650  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    7651  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    7652  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    7653  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    7654  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    7655  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    7656  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    7657  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    7658  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    7659  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    7660  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    7661  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    7662  : begin
              real_value= 32743;
              imag_value=1070;
            end
    7663  : begin
              real_value= 31843;
              imag_value=7699;
            end
    7664  : begin
              real_value= 29615;
              imag_value=14006;
            end
    7665  : begin
              real_value= 26152;
              imag_value=19729;
            end
    7666  : begin
              real_value= 21600;
              imag_value=24630;
            end
    7667  : begin
              real_value= 16148;
              imag_value=28506;
            end
    7668  : begin
              real_value= 10021;
              imag_value=31191;
            end
    7669  : begin
              real_value= 3476;
              imag_value=32575;
            end
    7670  : begin
              real_value= -3210;
              imag_value=32603;
            end
    7671  : begin
              real_value= -9765;
              imag_value=31271;
            end
    7672  : begin
              real_value= -15914;
              imag_value=28636;
            end
    7673  : begin
              real_value= -21399;
              imag_value=24806;
            end
    7674  : begin
              real_value= -25990;
              imag_value=19943;
            end
    7675  : begin
              real_value= -29499;
              imag_value=14248;
            end
    7676  : begin
              real_value= -31779;
              imag_value=7959;
            end
    7677  : begin
              real_value= -32733;
              imag_value=1338;
            end
    7678  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    7679  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    7680  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    7681  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    7682  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    7683  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    7684  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    7685  : begin
              real_value= 802;
              imag_value=-32750;
            end
    7686  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    7687  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    7688  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    7689  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    7690  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    7691  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    7692  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    7693  : begin
              real_value= 32629;
              imag_value=2942;
            end
    7694  : begin
              real_value= 31351;
              imag_value=9508;
            end
    7695  : begin
              real_value= 28766;
              imag_value=15678;
            end
    7696  : begin
              real_value= 24981;
              imag_value=21194;
            end
    7697  : begin
              real_value= 20154;
              imag_value=25826;
            end
    7698  : begin
              real_value= 14489;
              imag_value=29382;
            end
    7699  : begin
              real_value= 8219;
              imag_value=31713;
            end
    7700  : begin
              real_value= 1606;
              imag_value=32721;
            end
    7701  : begin
              real_value= -5071;
              imag_value=32365;
            end
    7702  : begin
              real_value= -11539;
              imag_value=30661;
            end
    7703  : begin
              real_value= -17525;
              imag_value=27678;
            end
    7704  : begin
              real_value= -22782;
              imag_value=23541;
            end
    7705  : begin
              real_value= -27090;
              imag_value=18423;
            end
    7706  : begin
              real_value= -30267;
              imag_value=12537;
            end
    7707  : begin
              real_value= -32183;
              imag_value=6127;
            end
    7708  : begin
              real_value= -32757;
              imag_value=-535;
            end
    7709  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    7710  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    7711  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    7712  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    7713  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    7714  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    7715  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    7716  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    7717  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    7718  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    7719  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    7720  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    7721  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    7722  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    7723  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    7724  : begin
              real_value= 32407;
              imag_value=4806;
            end
    7725  : begin
              real_value= 30755;
              imag_value=11289;
            end
    7726  : begin
              real_value= 27820;
              imag_value=17299;
            end
    7727  : begin
              real_value= 23726;
              imag_value=22589;
            end
    7728  : begin
              real_value= 18644;
              imag_value=26938;
            end
    7729  : begin
              real_value= 12784;
              imag_value=30163;
            end
    7730  : begin
              real_value= 6390;
              imag_value=32131;
            end
    7731  : begin
              real_value= -267;
              imag_value=32759;
            end
    7732  : begin
              real_value= -6915;
              imag_value=32022;
            end
    7733  : begin
              real_value= -13274;
              imag_value=29950;
            end
    7734  : begin
              real_value= -19081;
              imag_value=26630;
            end
    7735  : begin
              real_value= -24092;
              imag_value=22199;
            end
    7736  : begin
              real_value= -28100;
              imag_value=16842;
            end
    7737  : begin
              real_value= -30935;
              imag_value=10783;
            end
    7738  : begin
              real_value= -32481;
              imag_value=4275;
            end
    7739  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    7740  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    7741  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    7742  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    7743  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    7744  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    7745  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    7746  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    7747  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    7748  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    7749  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    7750  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    7751  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    7752  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    7753  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    7754  : begin
              real_value= 32760;
              imag_value=0;
            end
    7755  : begin
              real_value= 32077;
              imag_value=6654;
            end
    7756  : begin
              real_value= 30057;
              imag_value=13030;
            end
    7757  : begin
              real_value= 26784;
              imag_value=18863;
            end
    7758  : begin
              real_value= 22395;
              imag_value=23911;
            end
    7759  : begin
              real_value= 17072;
              imag_value=27961;
            end
    7760  : begin
              real_value= 11036;
              imag_value=30846;
            end
    7761  : begin
              real_value= 4540;
              imag_value=32445;
            end
    7762  : begin
              real_value= -2142;
              imag_value=32691;
            end
    7763  : begin
              real_value= -8737;
              imag_value=31575;
            end
    7764  : begin
              real_value= -14968;
              imag_value=29142;
            end
    7765  : begin
              real_value= -20575;
              imag_value=25494;
            end
    7766  : begin
              real_value= -25324;
              imag_value=20783;
            end
    7767  : begin
              real_value= -29017;
              imag_value=15206;
            end
    7768  : begin
              real_value= -31501;
              imag_value=8995;
            end
    7769  : begin
              real_value= -32673;
              imag_value=2408;
            end
    7770  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    7771  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    7772  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    7773  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    7774  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    7775  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    7776  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    7777  : begin
              real_value= -267;
              imag_value=-32759;
            end
    7778  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    7779  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    7780  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    7781  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    7782  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    7783  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    7784  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    7785  : begin
              real_value= 32707;
              imag_value=1874;
            end
    7786  : begin
              real_value= 31645;
              imag_value=8477;
            end
    7787  : begin
              real_value= 29263;
              imag_value=14728;
            end
    7788  : begin
              real_value= 25661;
              imag_value=20365;
            end
    7789  : begin
              real_value= 20988;
              imag_value=25154;
            end
    7790  : begin
              real_value= 15442;
              imag_value=28892;
            end
    7791  : begin
              real_value= 9253;
              imag_value=31426;
            end
    7792  : begin
              real_value= 2676;
              imag_value=32651;
            end
    7793  : begin
              real_value= -4009;
              imag_value=32515;
            end
    7794  : begin
              real_value= -10529;
              imag_value=31023;
            end
    7795  : begin
              real_value= -16611;
              imag_value=28236;
            end
    7796  : begin
              real_value= -22001;
              imag_value=24274;
            end
    7797  : begin
              real_value= -26472;
              imag_value=19299;
            end
    7798  : begin
              real_value= -29841;
              imag_value=13520;
            end
    7799  : begin
              real_value= -31965;
              imag_value=7177;
            end
    7800  : begin
              real_value= -32757;
              imag_value=535;
            end
    7801  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    7802  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    7803  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    7804  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    7805  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    7806  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    7807  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    7808  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    7809  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    7810  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    7811  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    7812  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    7813  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    7814  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    7815  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    7816  : begin
              real_value= 32547;
              imag_value=3742;
            end
    7817  : begin
              real_value= 31107;
              imag_value=10275;
            end
    7818  : begin
              real_value= 28371;
              imag_value=16380;
            end
    7819  : begin
              real_value= 24453;
              imag_value=21801;
            end
    7820  : begin
              real_value= 19515;
              imag_value=26314;
            end
    7821  : begin
              real_value= 13764;
              imag_value=29729;
            end
    7822  : begin
              real_value= 7438;
              imag_value=31905;
            end
    7823  : begin
              real_value= 802;
              imag_value=32750;
            end
    7824  : begin
              real_value= -5864;
              imag_value=32231;
            end
    7825  : begin
              real_value= -12288;
              imag_value=30369;
            end
    7826  : begin
              real_value= -18200;
              imag_value=27240;
            end
    7827  : begin
              real_value= -23354;
              imag_value=22974;
            end
    7828  : begin
              real_value= -27534;
              imag_value=17752;
            end
    7829  : begin
              real_value= -30565;
              imag_value=11790;
            end
    7830  : begin
              real_value= -32323;
              imag_value=5336;
            end
    7831  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    7832  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    7833  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    7834  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    7835  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    7836  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    7837  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    7838  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    7839  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    7840  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    7841  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    7842  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    7843  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    7844  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    7845  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    7846  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    7847  : begin
              real_value= 32278;
              imag_value=5599;
            end
    7848  : begin
              real_value= 30468;
              imag_value=12039;
            end
    7849  : begin
              real_value= 27387;
              imag_value=17977;
            end
    7850  : begin
              real_value= 23165;
              imag_value=23165;
            end
    7851  : begin
              real_value= 17977;
              imag_value=27387;
            end
    7852  : begin
              real_value= 12039;
              imag_value=30468;
            end
    7853  : begin
              real_value= 5599;
              imag_value=32278;
            end
    7854  : begin
              real_value= -1070;
              imag_value=32743;
            end
    7855  : begin
              real_value= -7699;
              imag_value=31843;
            end
    7856  : begin
              real_value= -14006;
              imag_value=29615;
            end
    7857  : begin
              real_value= -19729;
              imag_value=26152;
            end
    7858  : begin
              real_value= -24630;
              imag_value=21600;
            end
    7859  : begin
              real_value= -28506;
              imag_value=16148;
            end
    7860  : begin
              real_value= -31191;
              imag_value=10021;
            end
    7861  : begin
              real_value= -32575;
              imag_value=3476;
            end
    7862  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    7863  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    7864  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    7865  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    7866  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    7867  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    7868  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    7869  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    7870  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    7871  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    7872  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    7873  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    7874  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    7875  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    7876  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    7877  : begin
              real_value= 32750;
              imag_value=802;
            end
    7878  : begin
              real_value= 31905;
              imag_value=7438;
            end
    7879  : begin
              real_value= 29729;
              imag_value=13764;
            end
    7880  : begin
              real_value= 26314;
              imag_value=19515;
            end
    7881  : begin
              real_value= 21801;
              imag_value=24453;
            end
    7882  : begin
              real_value= 16380;
              imag_value=28371;
            end
    7883  : begin
              real_value= 10275;
              imag_value=31107;
            end
    7884  : begin
              real_value= 3742;
              imag_value=32547;
            end
    7885  : begin
              real_value= -2942;
              imag_value=32629;
            end
    7886  : begin
              real_value= -9508;
              imag_value=31351;
            end
    7887  : begin
              real_value= -15678;
              imag_value=28766;
            end
    7888  : begin
              real_value= -21194;
              imag_value=24981;
            end
    7889  : begin
              real_value= -25826;
              imag_value=20154;
            end
    7890  : begin
              real_value= -29382;
              imag_value=14489;
            end
    7891  : begin
              real_value= -31713;
              imag_value=8219;
            end
    7892  : begin
              real_value= -32721;
              imag_value=1606;
            end
    7893  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    7894  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    7895  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    7896  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    7897  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    7898  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    7899  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    7900  : begin
              real_value= 535;
              imag_value=-32757;
            end
    7901  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    7902  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    7903  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    7904  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    7905  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    7906  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    7907  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    7908  : begin
              real_value= 32651;
              imag_value=2676;
            end
    7909  : begin
              real_value= 31426;
              imag_value=9253;
            end
    7910  : begin
              real_value= 28892;
              imag_value=15442;
            end
    7911  : begin
              real_value= 25154;
              imag_value=20988;
            end
    7912  : begin
              real_value= 20365;
              imag_value=25661;
            end
    7913  : begin
              real_value= 14728;
              imag_value=29263;
            end
    7914  : begin
              real_value= 8477;
              imag_value=31645;
            end
    7915  : begin
              real_value= 1874;
              imag_value=32707;
            end
    7916  : begin
              real_value= -4806;
              imag_value=32407;
            end
    7917  : begin
              real_value= -11289;
              imag_value=30755;
            end
    7918  : begin
              real_value= -17299;
              imag_value=27820;
            end
    7919  : begin
              real_value= -22589;
              imag_value=23726;
            end
    7920  : begin
              real_value= -26938;
              imag_value=18644;
            end
    7921  : begin
              real_value= -30163;
              imag_value=12784;
            end
    7922  : begin
              real_value= -32131;
              imag_value=6390;
            end
    7923  : begin
              real_value= -32759;
              imag_value=-267;
            end
    7924  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    7925  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    7926  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    7927  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    7928  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    7929  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    7930  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    7931  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    7932  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    7933  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    7934  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    7935  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    7936  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    7937  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    7938  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    7939  : begin
              real_value= 32445;
              imag_value=4540;
            end
    7940  : begin
              real_value= 30846;
              imag_value=11036;
            end
    7941  : begin
              real_value= 27961;
              imag_value=17072;
            end
    7942  : begin
              real_value= 23911;
              imag_value=22395;
            end
    7943  : begin
              real_value= 18863;
              imag_value=26784;
            end
    7944  : begin
              real_value= 13030;
              imag_value=30057;
            end
    7945  : begin
              real_value= 6654;
              imag_value=32077;
            end
    7946  : begin
              real_value= 0;
              imag_value=32760;
            end
    7947  : begin
              real_value= -6654;
              imag_value=32077;
            end
    7948  : begin
              real_value= -13030;
              imag_value=30057;
            end
    7949  : begin
              real_value= -18863;
              imag_value=26784;
            end
    7950  : begin
              real_value= -23911;
              imag_value=22395;
            end
    7951  : begin
              real_value= -27961;
              imag_value=17072;
            end
    7952  : begin
              real_value= -30846;
              imag_value=11036;
            end
    7953  : begin
              real_value= -32445;
              imag_value=4540;
            end
    7954  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    7955  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    7956  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    7957  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    7958  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    7959  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    7960  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    7961  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    7962  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    7963  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    7964  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    7965  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    7966  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    7967  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    7968  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    7969  : begin
              real_value= 32759;
              imag_value=-267;
            end
    7970  : begin
              real_value= 32131;
              imag_value=6390;
            end
    7971  : begin
              real_value= 30163;
              imag_value=12784;
            end
    7972  : begin
              real_value= 26938;
              imag_value=18644;
            end
    7973  : begin
              real_value= 22589;
              imag_value=23726;
            end
    7974  : begin
              real_value= 17299;
              imag_value=27820;
            end
    7975  : begin
              real_value= 11289;
              imag_value=30755;
            end
    7976  : begin
              real_value= 4806;
              imag_value=32407;
            end
    7977  : begin
              real_value= -1874;
              imag_value=32707;
            end
    7978  : begin
              real_value= -8477;
              imag_value=31645;
            end
    7979  : begin
              real_value= -14728;
              imag_value=29263;
            end
    7980  : begin
              real_value= -20365;
              imag_value=25661;
            end
    7981  : begin
              real_value= -25154;
              imag_value=20988;
            end
    7982  : begin
              real_value= -28892;
              imag_value=15442;
            end
    7983  : begin
              real_value= -31426;
              imag_value=9253;
            end
    7984  : begin
              real_value= -32651;
              imag_value=2676;
            end
    7985  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    7986  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    7987  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    7988  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    7989  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    7990  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    7991  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    7992  : begin
              real_value= -535;
              imag_value=-32757;
            end
    7993  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    7994  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    7995  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    7996  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    7997  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    7998  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    7999  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    8000  : begin
              real_value= 32721;
              imag_value=1606;
            end
    8001  : begin
              real_value= 31713;
              imag_value=8219;
            end
    8002  : begin
              real_value= 29382;
              imag_value=14489;
            end
    8003  : begin
              real_value= 25826;
              imag_value=20154;
            end
    8004  : begin
              real_value= 21194;
              imag_value=24981;
            end
    8005  : begin
              real_value= 15678;
              imag_value=28766;
            end
    8006  : begin
              real_value= 9508;
              imag_value=31351;
            end
    8007  : begin
              real_value= 2942;
              imag_value=32629;
            end
    8008  : begin
              real_value= -3742;
              imag_value=32547;
            end
    8009  : begin
              real_value= -10275;
              imag_value=31107;
            end
    8010  : begin
              real_value= -16380;
              imag_value=28371;
            end
    8011  : begin
              real_value= -21801;
              imag_value=24453;
            end
    8012  : begin
              real_value= -26314;
              imag_value=19515;
            end
    8013  : begin
              real_value= -29729;
              imag_value=13764;
            end
    8014  : begin
              real_value= -31905;
              imag_value=7438;
            end
    8015  : begin
              real_value= -32750;
              imag_value=802;
            end
    8016  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    8017  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    8018  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    8019  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    8020  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    8021  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    8022  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    8023  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    8024  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    8025  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    8026  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    8027  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    8028  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    8029  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    8030  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    8031  : begin
              real_value= 32575;
              imag_value=3476;
            end
    8032  : begin
              real_value= 31191;
              imag_value=10021;
            end
    8033  : begin
              real_value= 28506;
              imag_value=16148;
            end
    8034  : begin
              real_value= 24630;
              imag_value=21600;
            end
    8035  : begin
              real_value= 19729;
              imag_value=26152;
            end
    8036  : begin
              real_value= 14006;
              imag_value=29615;
            end
    8037  : begin
              real_value= 7699;
              imag_value=31843;
            end
    8038  : begin
              real_value= 1070;
              imag_value=32743;
            end
    8039  : begin
              real_value= -5599;
              imag_value=32278;
            end
    8040  : begin
              real_value= -12039;
              imag_value=30468;
            end
    8041  : begin
              real_value= -17977;
              imag_value=27387;
            end
    8042  : begin
              real_value= -23165;
              imag_value=23165;
            end
    8043  : begin
              real_value= -27387;
              imag_value=17977;
            end
    8044  : begin
              real_value= -30468;
              imag_value=12039;
            end
    8045  : begin
              real_value= -32278;
              imag_value=5599;
            end
    8046  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    8047  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    8048  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    8049  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    8050  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    8051  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    8052  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    8053  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    8054  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    8055  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    8056  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    8057  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    8058  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    8059  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    8060  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    8061  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    8062  : begin
              real_value= 32323;
              imag_value=5336;
            end
    8063  : begin
              real_value= 30565;
              imag_value=11790;
            end
    8064  : begin
              real_value= 27534;
              imag_value=17752;
            end
    8065  : begin
              real_value= 23354;
              imag_value=22974;
            end
    8066  : begin
              real_value= 18200;
              imag_value=27240;
            end
    8067  : begin
              real_value= 12288;
              imag_value=30369;
            end
    8068  : begin
              real_value= 5864;
              imag_value=32231;
            end
    8069  : begin
              real_value= -802;
              imag_value=32750;
            end
    8070  : begin
              real_value= -7438;
              imag_value=31905;
            end
    8071  : begin
              real_value= -13764;
              imag_value=29729;
            end
    8072  : begin
              real_value= -19515;
              imag_value=26314;
            end
    8073  : begin
              real_value= -24453;
              imag_value=21801;
            end
    8074  : begin
              real_value= -28371;
              imag_value=16380;
            end
    8075  : begin
              real_value= -31107;
              imag_value=10275;
            end
    8076  : begin
              real_value= -32547;
              imag_value=3742;
            end
    8077  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    8078  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    8079  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    8080  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    8081  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    8082  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    8083  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    8084  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    8085  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    8086  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    8087  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    8088  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    8089  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    8090  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    8091  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    8092  : begin
              real_value= 32757;
              imag_value=535;
            end
    8093  : begin
              real_value= 31965;
              imag_value=7177;
            end
    8094  : begin
              real_value= 29841;
              imag_value=13520;
            end
    8095  : begin
              real_value= 26472;
              imag_value=19299;
            end
    8096  : begin
              real_value= 22001;
              imag_value=24274;
            end
    8097  : begin
              real_value= 16611;
              imag_value=28236;
            end
    8098  : begin
              real_value= 10529;
              imag_value=31023;
            end
    8099  : begin
              real_value= 4009;
              imag_value=32515;
            end
    8100  : begin
              real_value= -2676;
              imag_value=32651;
            end
    8101  : begin
              real_value= -9253;
              imag_value=31426;
            end
    8102  : begin
              real_value= -15442;
              imag_value=28892;
            end
    8103  : begin
              real_value= -20988;
              imag_value=25154;
            end
    8104  : begin
              real_value= -25661;
              imag_value=20365;
            end
    8105  : begin
              real_value= -29263;
              imag_value=14728;
            end
    8106  : begin
              real_value= -31645;
              imag_value=8477;
            end
    8107  : begin
              real_value= -32707;
              imag_value=1874;
            end
    8108  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    8109  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    8110  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    8111  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    8112  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    8113  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    8114  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    8115  : begin
              real_value= 267;
              imag_value=-32759;
            end
    8116  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    8117  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    8118  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    8119  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    8120  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    8121  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    8122  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    8123  : begin
              real_value= 32673;
              imag_value=2408;
            end
    8124  : begin
              real_value= 31501;
              imag_value=8995;
            end
    8125  : begin
              real_value= 29017;
              imag_value=15206;
            end
    8126  : begin
              real_value= 25324;
              imag_value=20783;
            end
    8127  : begin
              real_value= 20575;
              imag_value=25494;
            end
    8128  : begin
              real_value= 14968;
              imag_value=29142;
            end
    8129  : begin
              real_value= 8737;
              imag_value=31575;
            end
    8130  : begin
              real_value= 2142;
              imag_value=32691;
            end
    8131  : begin
              real_value= -4540;
              imag_value=32445;
            end
    8132  : begin
              real_value= -11036;
              imag_value=30846;
            end
    8133  : begin
              real_value= -17072;
              imag_value=27961;
            end
    8134  : begin
              real_value= -22395;
              imag_value=23911;
            end
    8135  : begin
              real_value= -26784;
              imag_value=18863;
            end
    8136  : begin
              real_value= -30057;
              imag_value=13030;
            end
    8137  : begin
              real_value= -32077;
              imag_value=6654;
            end
    8138  : begin
              real_value= -32760;
              imag_value=0;
            end
    8139  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    8140  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    8141  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    8142  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    8143  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    8144  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    8145  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    8146  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    8147  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    8148  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    8149  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    8150  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    8151  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    8152  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    8153  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    8154  : begin
              real_value= 32481;
              imag_value=4275;
            end
    8155  : begin
              real_value= 30935;
              imag_value=10783;
            end
    8156  : begin
              real_value= 28100;
              imag_value=16842;
            end
    8157  : begin
              real_value= 24092;
              imag_value=22199;
            end
    8158  : begin
              real_value= 19081;
              imag_value=26630;
            end
    8159  : begin
              real_value= 13274;
              imag_value=29950;
            end
    8160  : begin
              real_value= 6915;
              imag_value=32022;
            end
    8161  : begin
              real_value= 267;
              imag_value=32759;
            end
    8162  : begin
              real_value= -6390;
              imag_value=32131;
            end
    8163  : begin
              real_value= -12784;
              imag_value=30163;
            end
    8164  : begin
              real_value= -18644;
              imag_value=26938;
            end
    8165  : begin
              real_value= -23726;
              imag_value=22589;
            end
    8166  : begin
              real_value= -27820;
              imag_value=17299;
            end
    8167  : begin
              real_value= -30755;
              imag_value=11289;
            end
    8168  : begin
              real_value= -32407;
              imag_value=4806;
            end
    8169  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    8170  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    8171  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    8172  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    8173  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    8174  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    8175  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    8176  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    8177  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    8178  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    8179  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    8180  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    8181  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    8182  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    8183  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    8184  : begin
              real_value= 32757;
              imag_value=-535;
            end
    8185  : begin
              real_value= 32183;
              imag_value=6127;
            end
    8186  : begin
              real_value= 30267;
              imag_value=12537;
            end
    8187  : begin
              real_value= 27090;
              imag_value=18423;
            end
    8188  : begin
              real_value= 22782;
              imag_value=23541;
            end
    8189  : begin
              real_value= 17525;
              imag_value=27678;
            end
    8190  : begin
              real_value= 11539;
              imag_value=30661;
            end
    8191  : begin
              real_value= 5071;
              imag_value=32365;
            end
    8192  : begin
              real_value= -1606;
              imag_value=32721;
            end
    8193  : begin
              real_value= -8219;
              imag_value=31713;
            end
    8194  : begin
              real_value= -14489;
              imag_value=29382;
            end
    8195  : begin
              real_value= -20154;
              imag_value=25826;
            end
    8196  : begin
              real_value= -24981;
              imag_value=21194;
            end
    8197  : begin
              real_value= -28766;
              imag_value=15678;
            end
    8198  : begin
              real_value= -31351;
              imag_value=9508;
            end
    8199  : begin
              real_value= -32629;
              imag_value=2942;
            end
    8200  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    8201  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    8202  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    8203  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    8204  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    8205  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    8206  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    8207  : begin
              real_value= -802;
              imag_value=-32750;
            end
    8208  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    8209  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    8210  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    8211  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    8212  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    8213  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    8214  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    8215  : begin
              real_value= 32733;
              imag_value=1338;
            end
    8216  : begin
              real_value= 31779;
              imag_value=7959;
            end
    8217  : begin
              real_value= 29499;
              imag_value=14248;
            end
    8218  : begin
              real_value= 25990;
              imag_value=19943;
            end
    8219  : begin
              real_value= 21399;
              imag_value=24806;
            end
    8220  : begin
              real_value= 15914;
              imag_value=28636;
            end
    8221  : begin
              real_value= 9765;
              imag_value=31271;
            end
    8222  : begin
              real_value= 3210;
              imag_value=32603;
            end
    8223  : begin
              real_value= -3476;
              imag_value=32575;
            end
    8224  : begin
              real_value= -10021;
              imag_value=31191;
            end
    8225  : begin
              real_value= -16148;
              imag_value=28506;
            end
    8226  : begin
              real_value= -21600;
              imag_value=24630;
            end
    8227  : begin
              real_value= -26152;
              imag_value=19729;
            end
    8228  : begin
              real_value= -29615;
              imag_value=14006;
            end
    8229  : begin
              real_value= -31843;
              imag_value=7699;
            end
    8230  : begin
              real_value= -32743;
              imag_value=1070;
            end
    8231  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    8232  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    8233  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    8234  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    8235  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    8236  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    8237  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    8238  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    8239  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    8240  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    8241  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    8242  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    8243  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    8244  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    8245  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    8246  : begin
              real_value= 32603;
              imag_value=3210;
            end
    8247  : begin
              real_value= 31271;
              imag_value=9765;
            end
    8248  : begin
              real_value= 28636;
              imag_value=15914;
            end
    8249  : begin
              real_value= 24806;
              imag_value=21399;
            end
    8250  : begin
              real_value= 19943;
              imag_value=25990;
            end
    8251  : begin
              real_value= 14248;
              imag_value=29499;
            end
    8252  : begin
              real_value= 7959;
              imag_value=31779;
            end
    8253  : begin
              real_value= 1338;
              imag_value=32733;
            end
    8254  : begin
              real_value= -5336;
              imag_value=32323;
            end
    8255  : begin
              real_value= -11790;
              imag_value=30565;
            end
    8256  : begin
              real_value= -17752;
              imag_value=27534;
            end
    8257  : begin
              real_value= -22974;
              imag_value=23354;
            end
    8258  : begin
              real_value= -27240;
              imag_value=18200;
            end
    8259  : begin
              real_value= -30369;
              imag_value=12288;
            end
    8260  : begin
              real_value= -32231;
              imag_value=5864;
            end
    8261  : begin
              real_value= -32750;
              imag_value=-802;
            end
    8262  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    8263  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    8264  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    8265  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    8266  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    8267  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    8268  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    8269  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    8270  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    8271  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    8272  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    8273  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    8274  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    8275  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    8276  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    8277  : begin
              real_value= 32365;
              imag_value=5071;
            end
    8278  : begin
              real_value= 30661;
              imag_value=11539;
            end
    8279  : begin
              real_value= 27678;
              imag_value=17525;
            end
    8280  : begin
              real_value= 23541;
              imag_value=22782;
            end
    8281  : begin
              real_value= 18423;
              imag_value=27090;
            end
    8282  : begin
              real_value= 12537;
              imag_value=30267;
            end
    8283  : begin
              real_value= 6127;
              imag_value=32183;
            end
    8284  : begin
              real_value= -535;
              imag_value=32757;
            end
    8285  : begin
              real_value= -7177;
              imag_value=31965;
            end
    8286  : begin
              real_value= -13520;
              imag_value=29841;
            end
    8287  : begin
              real_value= -19299;
              imag_value=26472;
            end
    8288  : begin
              real_value= -24274;
              imag_value=22001;
            end
    8289  : begin
              real_value= -28236;
              imag_value=16611;
            end
    8290  : begin
              real_value= -31023;
              imag_value=10529;
            end
    8291  : begin
              real_value= -32515;
              imag_value=4009;
            end
    8292  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    8293  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    8294  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    8295  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    8296  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    8297  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    8298  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    8299  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    8300  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    8301  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    8302  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    8303  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    8304  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    8305  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    8306  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    8307  : begin
              real_value= 32759;
              imag_value=267;
            end
    8308  : begin
              real_value= 32022;
              imag_value=6915;
            end
    8309  : begin
              real_value= 29950;
              imag_value=13274;
            end
    8310  : begin
              real_value= 26630;
              imag_value=19081;
            end
    8311  : begin
              real_value= 22199;
              imag_value=24092;
            end
    8312  : begin
              real_value= 16842;
              imag_value=28100;
            end
    8313  : begin
              real_value= 10783;
              imag_value=30935;
            end
    8314  : begin
              real_value= 4275;
              imag_value=32481;
            end
    8315  : begin
              real_value= -2408;
              imag_value=32673;
            end
    8316  : begin
              real_value= -8995;
              imag_value=31501;
            end
    8317  : begin
              real_value= -15206;
              imag_value=29017;
            end
    8318  : begin
              real_value= -20783;
              imag_value=25324;
            end
    8319  : begin
              real_value= -25494;
              imag_value=20575;
            end
    8320  : begin
              real_value= -29142;
              imag_value=14968;
            end
    8321  : begin
              real_value= -31575;
              imag_value=8737;
            end
    8322  : begin
              real_value= -32691;
              imag_value=2142;
            end
    8323  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    8324  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    8325  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    8326  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    8327  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    8328  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    8329  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    8330  : begin
              real_value= 0;
              imag_value=-32760;
            end
    8331  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    8332  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    8333  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    8334  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    8335  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    8336  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    8337  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    8338  : begin
              real_value= 32691;
              imag_value=2142;
            end
    8339  : begin
              real_value= 31575;
              imag_value=8737;
            end
    8340  : begin
              real_value= 29142;
              imag_value=14968;
            end
    8341  : begin
              real_value= 25494;
              imag_value=20575;
            end
    8342  : begin
              real_value= 20783;
              imag_value=25324;
            end
    8343  : begin
              real_value= 15206;
              imag_value=29017;
            end
    8344  : begin
              real_value= 8995;
              imag_value=31501;
            end
    8345  : begin
              real_value= 2408;
              imag_value=32673;
            end
    8346  : begin
              real_value= -4275;
              imag_value=32481;
            end
    8347  : begin
              real_value= -10783;
              imag_value=30935;
            end
    8348  : begin
              real_value= -16842;
              imag_value=28100;
            end
    8349  : begin
              real_value= -22199;
              imag_value=24092;
            end
    8350  : begin
              real_value= -26630;
              imag_value=19081;
            end
    8351  : begin
              real_value= -29950;
              imag_value=13274;
            end
    8352  : begin
              real_value= -32022;
              imag_value=6915;
            end
    8353  : begin
              real_value= -32759;
              imag_value=267;
            end
    8354  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    8355  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    8356  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    8357  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    8358  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    8359  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    8360  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    8361  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    8362  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    8363  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    8364  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    8365  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    8366  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    8367  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    8368  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    8369  : begin
              real_value= 32515;
              imag_value=4009;
            end
    8370  : begin
              real_value= 31023;
              imag_value=10529;
            end
    8371  : begin
              real_value= 28236;
              imag_value=16611;
            end
    8372  : begin
              real_value= 24274;
              imag_value=22001;
            end
    8373  : begin
              real_value= 19299;
              imag_value=26472;
            end
    8374  : begin
              real_value= 13520;
              imag_value=29841;
            end
    8375  : begin
              real_value= 7177;
              imag_value=31965;
            end
    8376  : begin
              real_value= 535;
              imag_value=32757;
            end
    8377  : begin
              real_value= -6127;
              imag_value=32183;
            end
    8378  : begin
              real_value= -12537;
              imag_value=30267;
            end
    8379  : begin
              real_value= -18423;
              imag_value=27090;
            end
    8380  : begin
              real_value= -23541;
              imag_value=22782;
            end
    8381  : begin
              real_value= -27678;
              imag_value=17525;
            end
    8382  : begin
              real_value= -30661;
              imag_value=11539;
            end
    8383  : begin
              real_value= -32365;
              imag_value=5071;
            end
    8384  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    8385  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    8386  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    8387  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    8388  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    8389  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    8390  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    8391  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    8392  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    8393  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    8394  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    8395  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    8396  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    8397  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    8398  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    8399  : begin
              real_value= 32750;
              imag_value=-802;
            end
    8400  : begin
              real_value= 32231;
              imag_value=5864;
            end
    8401  : begin
              real_value= 30369;
              imag_value=12288;
            end
    8402  : begin
              real_value= 27240;
              imag_value=18200;
            end
    8403  : begin
              real_value= 22974;
              imag_value=23354;
            end
    8404  : begin
              real_value= 17752;
              imag_value=27534;
            end
    8405  : begin
              real_value= 11790;
              imag_value=30565;
            end
    8406  : begin
              real_value= 5336;
              imag_value=32323;
            end
    8407  : begin
              real_value= -1338;
              imag_value=32733;
            end
    8408  : begin
              real_value= -7959;
              imag_value=31779;
            end
    8409  : begin
              real_value= -14248;
              imag_value=29499;
            end
    8410  : begin
              real_value= -19943;
              imag_value=25990;
            end
    8411  : begin
              real_value= -24806;
              imag_value=21399;
            end
    8412  : begin
              real_value= -28636;
              imag_value=15914;
            end
    8413  : begin
              real_value= -31271;
              imag_value=9765;
            end
    8414  : begin
              real_value= -32603;
              imag_value=3210;
            end
    8415  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    8416  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    8417  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    8418  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    8419  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    8420  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    8421  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    8422  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    8423  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    8424  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    8425  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    8426  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    8427  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    8428  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    8429  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    8430  : begin
              real_value= 32743;
              imag_value=1070;
            end
    8431  : begin
              real_value= 31843;
              imag_value=7699;
            end
    8432  : begin
              real_value= 29615;
              imag_value=14006;
            end
    8433  : begin
              real_value= 26152;
              imag_value=19729;
            end
    8434  : begin
              real_value= 21600;
              imag_value=24630;
            end
    8435  : begin
              real_value= 16148;
              imag_value=28506;
            end
    8436  : begin
              real_value= 10021;
              imag_value=31191;
            end
    8437  : begin
              real_value= 3476;
              imag_value=32575;
            end
    8438  : begin
              real_value= -3210;
              imag_value=32603;
            end
    8439  : begin
              real_value= -9765;
              imag_value=31271;
            end
    8440  : begin
              real_value= -15914;
              imag_value=28636;
            end
    8441  : begin
              real_value= -21399;
              imag_value=24806;
            end
    8442  : begin
              real_value= -25990;
              imag_value=19943;
            end
    8443  : begin
              real_value= -29499;
              imag_value=14248;
            end
    8444  : begin
              real_value= -31779;
              imag_value=7959;
            end
    8445  : begin
              real_value= -32733;
              imag_value=1338;
            end
    8446  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    8447  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    8448  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    8449  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    8450  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    8451  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    8452  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    8453  : begin
              real_value= 802;
              imag_value=-32750;
            end
    8454  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    8455  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    8456  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    8457  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    8458  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    8459  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    8460  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    8461  : begin
              real_value= 32629;
              imag_value=2942;
            end
    8462  : begin
              real_value= 31351;
              imag_value=9508;
            end
    8463  : begin
              real_value= 28766;
              imag_value=15678;
            end
    8464  : begin
              real_value= 24981;
              imag_value=21194;
            end
    8465  : begin
              real_value= 20154;
              imag_value=25826;
            end
    8466  : begin
              real_value= 14489;
              imag_value=29382;
            end
    8467  : begin
              real_value= 8219;
              imag_value=31713;
            end
    8468  : begin
              real_value= 1606;
              imag_value=32721;
            end
    8469  : begin
              real_value= -5071;
              imag_value=32365;
            end
    8470  : begin
              real_value= -11539;
              imag_value=30661;
            end
    8471  : begin
              real_value= -17525;
              imag_value=27678;
            end
    8472  : begin
              real_value= -22782;
              imag_value=23541;
            end
    8473  : begin
              real_value= -27090;
              imag_value=18423;
            end
    8474  : begin
              real_value= -30267;
              imag_value=12537;
            end
    8475  : begin
              real_value= -32183;
              imag_value=6127;
            end
    8476  : begin
              real_value= -32757;
              imag_value=-535;
            end
    8477  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    8478  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    8479  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    8480  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    8481  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    8482  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    8483  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    8484  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    8485  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    8486  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    8487  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    8488  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    8489  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    8490  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    8491  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    8492  : begin
              real_value= 32407;
              imag_value=4806;
            end
    8493  : begin
              real_value= 30755;
              imag_value=11289;
            end
    8494  : begin
              real_value= 27820;
              imag_value=17299;
            end
    8495  : begin
              real_value= 23726;
              imag_value=22589;
            end
    8496  : begin
              real_value= 18644;
              imag_value=26938;
            end
    8497  : begin
              real_value= 12784;
              imag_value=30163;
            end
    8498  : begin
              real_value= 6390;
              imag_value=32131;
            end
    8499  : begin
              real_value= -267;
              imag_value=32759;
            end
    8500  : begin
              real_value= -6915;
              imag_value=32022;
            end
    8501  : begin
              real_value= -13274;
              imag_value=29950;
            end
    8502  : begin
              real_value= -19081;
              imag_value=26630;
            end
    8503  : begin
              real_value= -24092;
              imag_value=22199;
            end
    8504  : begin
              real_value= -28100;
              imag_value=16842;
            end
    8505  : begin
              real_value= -30935;
              imag_value=10783;
            end
    8506  : begin
              real_value= -32481;
              imag_value=4275;
            end
    8507  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    8508  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    8509  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    8510  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    8511  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    8512  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    8513  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    8514  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    8515  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    8516  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    8517  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    8518  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    8519  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    8520  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    8521  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    8522  : begin
              real_value= 32760;
              imag_value=0;
            end
    8523  : begin
              real_value= 32077;
              imag_value=6654;
            end
    8524  : begin
              real_value= 30057;
              imag_value=13030;
            end
    8525  : begin
              real_value= 26784;
              imag_value=18863;
            end
    8526  : begin
              real_value= 22395;
              imag_value=23911;
            end
    8527  : begin
              real_value= 17072;
              imag_value=27961;
            end
    8528  : begin
              real_value= 11036;
              imag_value=30846;
            end
    8529  : begin
              real_value= 4540;
              imag_value=32445;
            end
    8530  : begin
              real_value= -2142;
              imag_value=32691;
            end
    8531  : begin
              real_value= -8737;
              imag_value=31575;
            end
    8532  : begin
              real_value= -14968;
              imag_value=29142;
            end
    8533  : begin
              real_value= -20575;
              imag_value=25494;
            end
    8534  : begin
              real_value= -25324;
              imag_value=20783;
            end
    8535  : begin
              real_value= -29017;
              imag_value=15206;
            end
    8536  : begin
              real_value= -31501;
              imag_value=8995;
            end
    8537  : begin
              real_value= -32673;
              imag_value=2408;
            end
    8538  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    8539  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    8540  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    8541  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    8542  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    8543  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    8544  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    8545  : begin
              real_value= -267;
              imag_value=-32759;
            end
    8546  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    8547  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    8548  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    8549  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    8550  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    8551  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    8552  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    8553  : begin
              real_value= 32707;
              imag_value=1874;
            end
    8554  : begin
              real_value= 31645;
              imag_value=8477;
            end
    8555  : begin
              real_value= 29263;
              imag_value=14728;
            end
    8556  : begin
              real_value= 25661;
              imag_value=20365;
            end
    8557  : begin
              real_value= 20988;
              imag_value=25154;
            end
    8558  : begin
              real_value= 15442;
              imag_value=28892;
            end
    8559  : begin
              real_value= 9253;
              imag_value=31426;
            end
    8560  : begin
              real_value= 2676;
              imag_value=32651;
            end
    8561  : begin
              real_value= -4009;
              imag_value=32515;
            end
    8562  : begin
              real_value= -10529;
              imag_value=31023;
            end
    8563  : begin
              real_value= -16611;
              imag_value=28236;
            end
    8564  : begin
              real_value= -22001;
              imag_value=24274;
            end
    8565  : begin
              real_value= -26472;
              imag_value=19299;
            end
    8566  : begin
              real_value= -29841;
              imag_value=13520;
            end
    8567  : begin
              real_value= -31965;
              imag_value=7177;
            end
    8568  : begin
              real_value= -32757;
              imag_value=535;
            end
    8569  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    8570  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    8571  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    8572  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    8573  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    8574  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    8575  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    8576  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    8577  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    8578  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    8579  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    8580  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    8581  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    8582  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    8583  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    8584  : begin
              real_value= 32547;
              imag_value=3742;
            end
    8585  : begin
              real_value= 31107;
              imag_value=10275;
            end
    8586  : begin
              real_value= 28371;
              imag_value=16380;
            end
    8587  : begin
              real_value= 24453;
              imag_value=21801;
            end
    8588  : begin
              real_value= 19515;
              imag_value=26314;
            end
    8589  : begin
              real_value= 13764;
              imag_value=29729;
            end
    8590  : begin
              real_value= 7438;
              imag_value=31905;
            end
    8591  : begin
              real_value= 802;
              imag_value=32750;
            end
    8592  : begin
              real_value= -5864;
              imag_value=32231;
            end
    8593  : begin
              real_value= -12288;
              imag_value=30369;
            end
    8594  : begin
              real_value= -18200;
              imag_value=27240;
            end
    8595  : begin
              real_value= -23354;
              imag_value=22974;
            end
    8596  : begin
              real_value= -27534;
              imag_value=17752;
            end
    8597  : begin
              real_value= -30565;
              imag_value=11790;
            end
    8598  : begin
              real_value= -32323;
              imag_value=5336;
            end
    8599  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    8600  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    8601  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    8602  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    8603  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    8604  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    8605  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    8606  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    8607  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    8608  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    8609  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    8610  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    8611  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    8612  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    8613  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    8614  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    8615  : begin
              real_value= 32278;
              imag_value=5599;
            end
    8616  : begin
              real_value= 30468;
              imag_value=12039;
            end
    8617  : begin
              real_value= 27387;
              imag_value=17977;
            end
    8618  : begin
              real_value= 23165;
              imag_value=23165;
            end
    8619  : begin
              real_value= 17977;
              imag_value=27387;
            end
    8620  : begin
              real_value= 12039;
              imag_value=30468;
            end
    8621  : begin
              real_value= 5599;
              imag_value=32278;
            end
    8622  : begin
              real_value= -1070;
              imag_value=32743;
            end
    8623  : begin
              real_value= -7699;
              imag_value=31843;
            end
    8624  : begin
              real_value= -14006;
              imag_value=29615;
            end
    8625  : begin
              real_value= -19729;
              imag_value=26152;
            end
    8626  : begin
              real_value= -24630;
              imag_value=21600;
            end
    8627  : begin
              real_value= -28506;
              imag_value=16148;
            end
    8628  : begin
              real_value= -31191;
              imag_value=10021;
            end
    8629  : begin
              real_value= -32575;
              imag_value=3476;
            end
    8630  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    8631  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    8632  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    8633  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    8634  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    8635  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    8636  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    8637  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    8638  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    8639  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    8640  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    8641  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    8642  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    8643  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    8644  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    8645  : begin
              real_value= 32750;
              imag_value=802;
            end
    8646  : begin
              real_value= 31905;
              imag_value=7438;
            end
    8647  : begin
              real_value= 29729;
              imag_value=13764;
            end
    8648  : begin
              real_value= 26314;
              imag_value=19515;
            end
    8649  : begin
              real_value= 21801;
              imag_value=24453;
            end
    8650  : begin
              real_value= 16380;
              imag_value=28371;
            end
    8651  : begin
              real_value= 10275;
              imag_value=31107;
            end
    8652  : begin
              real_value= 3742;
              imag_value=32547;
            end
    8653  : begin
              real_value= -2942;
              imag_value=32629;
            end
    8654  : begin
              real_value= -9508;
              imag_value=31351;
            end
    8655  : begin
              real_value= -15678;
              imag_value=28766;
            end
    8656  : begin
              real_value= -21194;
              imag_value=24981;
            end
    8657  : begin
              real_value= -25826;
              imag_value=20154;
            end
    8658  : begin
              real_value= -29382;
              imag_value=14489;
            end
    8659  : begin
              real_value= -31713;
              imag_value=8219;
            end
    8660  : begin
              real_value= -32721;
              imag_value=1606;
            end
    8661  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    8662  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    8663  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    8664  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    8665  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    8666  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    8667  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    8668  : begin
              real_value= 535;
              imag_value=-32757;
            end
    8669  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    8670  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    8671  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    8672  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    8673  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    8674  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    8675  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    8676  : begin
              real_value= 32651;
              imag_value=2676;
            end
    8677  : begin
              real_value= 31426;
              imag_value=9253;
            end
    8678  : begin
              real_value= 28892;
              imag_value=15442;
            end
    8679  : begin
              real_value= 25154;
              imag_value=20988;
            end
    8680  : begin
              real_value= 20365;
              imag_value=25661;
            end
    8681  : begin
              real_value= 14728;
              imag_value=29263;
            end
    8682  : begin
              real_value= 8477;
              imag_value=31645;
            end
    8683  : begin
              real_value= 1874;
              imag_value=32707;
            end
    8684  : begin
              real_value= -4806;
              imag_value=32407;
            end
    8685  : begin
              real_value= -11289;
              imag_value=30755;
            end
    8686  : begin
              real_value= -17299;
              imag_value=27820;
            end
    8687  : begin
              real_value= -22589;
              imag_value=23726;
            end
    8688  : begin
              real_value= -26938;
              imag_value=18644;
            end
    8689  : begin
              real_value= -30163;
              imag_value=12784;
            end
    8690  : begin
              real_value= -32131;
              imag_value=6390;
            end
    8691  : begin
              real_value= -32759;
              imag_value=-267;
            end
    8692  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    8693  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    8694  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    8695  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    8696  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    8697  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    8698  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    8699  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    8700  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    8701  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    8702  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    8703  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    8704  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    8705  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    8706  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    8707  : begin
              real_value= 32445;
              imag_value=4540;
            end
    8708  : begin
              real_value= 30846;
              imag_value=11036;
            end
    8709  : begin
              real_value= 27961;
              imag_value=17072;
            end
    8710  : begin
              real_value= 23911;
              imag_value=22395;
            end
    8711  : begin
              real_value= 18863;
              imag_value=26784;
            end
    8712  : begin
              real_value= 13030;
              imag_value=30057;
            end
    8713  : begin
              real_value= 6654;
              imag_value=32077;
            end
    8714  : begin
              real_value= 0;
              imag_value=32760;
            end
    8715  : begin
              real_value= -6654;
              imag_value=32077;
            end
    8716  : begin
              real_value= -13030;
              imag_value=30057;
            end
    8717  : begin
              real_value= -18863;
              imag_value=26784;
            end
    8718  : begin
              real_value= -23911;
              imag_value=22395;
            end
    8719  : begin
              real_value= -27961;
              imag_value=17072;
            end
    8720  : begin
              real_value= -30846;
              imag_value=11036;
            end
    8721  : begin
              real_value= -32445;
              imag_value=4540;
            end
    8722  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    8723  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    8724  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    8725  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    8726  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    8727  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    8728  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    8729  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    8730  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    8731  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    8732  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    8733  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    8734  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    8735  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    8736  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    8737  : begin
              real_value= 32759;
              imag_value=-267;
            end
    8738  : begin
              real_value= 32131;
              imag_value=6390;
            end
    8739  : begin
              real_value= 30163;
              imag_value=12784;
            end
    8740  : begin
              real_value= 26938;
              imag_value=18644;
            end
    8741  : begin
              real_value= 22589;
              imag_value=23726;
            end
    8742  : begin
              real_value= 17299;
              imag_value=27820;
            end
    8743  : begin
              real_value= 11289;
              imag_value=30755;
            end
    8744  : begin
              real_value= 4806;
              imag_value=32407;
            end
    8745  : begin
              real_value= -1874;
              imag_value=32707;
            end
    8746  : begin
              real_value= -8477;
              imag_value=31645;
            end
    8747  : begin
              real_value= -14728;
              imag_value=29263;
            end
    8748  : begin
              real_value= -20365;
              imag_value=25661;
            end
    8749  : begin
              real_value= -25154;
              imag_value=20988;
            end
    8750  : begin
              real_value= -28892;
              imag_value=15442;
            end
    8751  : begin
              real_value= -31426;
              imag_value=9253;
            end
    8752  : begin
              real_value= -32651;
              imag_value=2676;
            end
    8753  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    8754  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    8755  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    8756  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    8757  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    8758  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    8759  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    8760  : begin
              real_value= -535;
              imag_value=-32757;
            end
    8761  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    8762  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    8763  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    8764  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    8765  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    8766  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    8767  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    8768  : begin
              real_value= 32721;
              imag_value=1606;
            end
    8769  : begin
              real_value= 31713;
              imag_value=8219;
            end
    8770  : begin
              real_value= 29382;
              imag_value=14489;
            end
    8771  : begin
              real_value= 25826;
              imag_value=20154;
            end
    8772  : begin
              real_value= 21194;
              imag_value=24981;
            end
    8773  : begin
              real_value= 15678;
              imag_value=28766;
            end
    8774  : begin
              real_value= 9508;
              imag_value=31351;
            end
    8775  : begin
              real_value= 2942;
              imag_value=32629;
            end
    8776  : begin
              real_value= -3742;
              imag_value=32547;
            end
    8777  : begin
              real_value= -10275;
              imag_value=31107;
            end
    8778  : begin
              real_value= -16380;
              imag_value=28371;
            end
    8779  : begin
              real_value= -21801;
              imag_value=24453;
            end
    8780  : begin
              real_value= -26314;
              imag_value=19515;
            end
    8781  : begin
              real_value= -29729;
              imag_value=13764;
            end
    8782  : begin
              real_value= -31905;
              imag_value=7438;
            end
    8783  : begin
              real_value= -32750;
              imag_value=802;
            end
    8784  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    8785  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    8786  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    8787  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    8788  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    8789  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    8790  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    8791  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    8792  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    8793  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    8794  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    8795  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    8796  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    8797  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    8798  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    8799  : begin
              real_value= 32575;
              imag_value=3476;
            end
    8800  : begin
              real_value= 31191;
              imag_value=10021;
            end
    8801  : begin
              real_value= 28506;
              imag_value=16148;
            end
    8802  : begin
              real_value= 24630;
              imag_value=21600;
            end
    8803  : begin
              real_value= 19729;
              imag_value=26152;
            end
    8804  : begin
              real_value= 14006;
              imag_value=29615;
            end
    8805  : begin
              real_value= 7699;
              imag_value=31843;
            end
    8806  : begin
              real_value= 1070;
              imag_value=32743;
            end
    8807  : begin
              real_value= -5599;
              imag_value=32278;
            end
    8808  : begin
              real_value= -12039;
              imag_value=30468;
            end
    8809  : begin
              real_value= -17977;
              imag_value=27387;
            end
    8810  : begin
              real_value= -23165;
              imag_value=23165;
            end
    8811  : begin
              real_value= -27387;
              imag_value=17977;
            end
    8812  : begin
              real_value= -30468;
              imag_value=12039;
            end
    8813  : begin
              real_value= -32278;
              imag_value=5599;
            end
    8814  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    8815  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    8816  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    8817  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    8818  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    8819  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    8820  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    8821  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    8822  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    8823  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    8824  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    8825  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    8826  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    8827  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    8828  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    8829  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    8830  : begin
              real_value= 32323;
              imag_value=5336;
            end
    8831  : begin
              real_value= 30565;
              imag_value=11790;
            end
    8832  : begin
              real_value= 27534;
              imag_value=17752;
            end
    8833  : begin
              real_value= 23354;
              imag_value=22974;
            end
    8834  : begin
              real_value= 18200;
              imag_value=27240;
            end
    8835  : begin
              real_value= 12288;
              imag_value=30369;
            end
    8836  : begin
              real_value= 5864;
              imag_value=32231;
            end
    8837  : begin
              real_value= -802;
              imag_value=32750;
            end
    8838  : begin
              real_value= -7438;
              imag_value=31905;
            end
    8839  : begin
              real_value= -13764;
              imag_value=29729;
            end
    8840  : begin
              real_value= -19515;
              imag_value=26314;
            end
    8841  : begin
              real_value= -24453;
              imag_value=21801;
            end
    8842  : begin
              real_value= -28371;
              imag_value=16380;
            end
    8843  : begin
              real_value= -31107;
              imag_value=10275;
            end
    8844  : begin
              real_value= -32547;
              imag_value=3742;
            end
    8845  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    8846  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    8847  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    8848  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    8849  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    8850  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    8851  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    8852  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    8853  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    8854  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    8855  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    8856  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    8857  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    8858  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    8859  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    8860  : begin
              real_value= 32757;
              imag_value=535;
            end
    8861  : begin
              real_value= 31965;
              imag_value=7177;
            end
    8862  : begin
              real_value= 29841;
              imag_value=13520;
            end
    8863  : begin
              real_value= 26472;
              imag_value=19299;
            end
    8864  : begin
              real_value= 22001;
              imag_value=24274;
            end
    8865  : begin
              real_value= 16611;
              imag_value=28236;
            end
    8866  : begin
              real_value= 10529;
              imag_value=31023;
            end
    8867  : begin
              real_value= 4009;
              imag_value=32515;
            end
    8868  : begin
              real_value= -2676;
              imag_value=32651;
            end
    8869  : begin
              real_value= -9253;
              imag_value=31426;
            end
    8870  : begin
              real_value= -15442;
              imag_value=28892;
            end
    8871  : begin
              real_value= -20988;
              imag_value=25154;
            end
    8872  : begin
              real_value= -25661;
              imag_value=20365;
            end
    8873  : begin
              real_value= -29263;
              imag_value=14728;
            end
    8874  : begin
              real_value= -31645;
              imag_value=8477;
            end
    8875  : begin
              real_value= -32707;
              imag_value=1874;
            end
    8876  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    8877  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    8878  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    8879  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    8880  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    8881  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    8882  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    8883  : begin
              real_value= 267;
              imag_value=-32759;
            end
    8884  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    8885  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    8886  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    8887  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    8888  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    8889  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    8890  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    8891  : begin
              real_value= 32673;
              imag_value=2408;
            end
    8892  : begin
              real_value= 31501;
              imag_value=8995;
            end
    8893  : begin
              real_value= 29017;
              imag_value=15206;
            end
    8894  : begin
              real_value= 25324;
              imag_value=20783;
            end
    8895  : begin
              real_value= 20575;
              imag_value=25494;
            end
    8896  : begin
              real_value= 14968;
              imag_value=29142;
            end
    8897  : begin
              real_value= 8737;
              imag_value=31575;
            end
    8898  : begin
              real_value= 2142;
              imag_value=32691;
            end
    8899  : begin
              real_value= -4540;
              imag_value=32445;
            end
    8900  : begin
              real_value= -11036;
              imag_value=30846;
            end
    8901  : begin
              real_value= -17072;
              imag_value=27961;
            end
    8902  : begin
              real_value= -22395;
              imag_value=23911;
            end
    8903  : begin
              real_value= -26784;
              imag_value=18863;
            end
    8904  : begin
              real_value= -30057;
              imag_value=13030;
            end
    8905  : begin
              real_value= -32077;
              imag_value=6654;
            end
    8906  : begin
              real_value= -32760;
              imag_value=0;
            end
    8907  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    8908  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    8909  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    8910  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    8911  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    8912  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    8913  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    8914  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    8915  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    8916  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    8917  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    8918  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    8919  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    8920  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    8921  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    8922  : begin
              real_value= 32481;
              imag_value=4275;
            end
    8923  : begin
              real_value= 30935;
              imag_value=10783;
            end
    8924  : begin
              real_value= 28100;
              imag_value=16842;
            end
    8925  : begin
              real_value= 24092;
              imag_value=22199;
            end
    8926  : begin
              real_value= 19081;
              imag_value=26630;
            end
    8927  : begin
              real_value= 13274;
              imag_value=29950;
            end
    8928  : begin
              real_value= 6915;
              imag_value=32022;
            end
    8929  : begin
              real_value= 267;
              imag_value=32759;
            end
    8930  : begin
              real_value= -6390;
              imag_value=32131;
            end
    8931  : begin
              real_value= -12784;
              imag_value=30163;
            end
    8932  : begin
              real_value= -18644;
              imag_value=26938;
            end
    8933  : begin
              real_value= -23726;
              imag_value=22589;
            end
    8934  : begin
              real_value= -27820;
              imag_value=17299;
            end
    8935  : begin
              real_value= -30755;
              imag_value=11289;
            end
    8936  : begin
              real_value= -32407;
              imag_value=4806;
            end
    8937  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    8938  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    8939  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    8940  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    8941  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    8942  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    8943  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    8944  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    8945  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    8946  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    8947  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    8948  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    8949  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    8950  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    8951  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    8952  : begin
              real_value= 32757;
              imag_value=-535;
            end
    8953  : begin
              real_value= 32183;
              imag_value=6127;
            end
    8954  : begin
              real_value= 30267;
              imag_value=12537;
            end
    8955  : begin
              real_value= 27090;
              imag_value=18423;
            end
    8956  : begin
              real_value= 22782;
              imag_value=23541;
            end
    8957  : begin
              real_value= 17525;
              imag_value=27678;
            end
    8958  : begin
              real_value= 11539;
              imag_value=30661;
            end
    8959  : begin
              real_value= 5071;
              imag_value=32365;
            end
    8960  : begin
              real_value= -1606;
              imag_value=32721;
            end
    8961  : begin
              real_value= -8219;
              imag_value=31713;
            end
    8962  : begin
              real_value= -14489;
              imag_value=29382;
            end
    8963  : begin
              real_value= -20154;
              imag_value=25826;
            end
    8964  : begin
              real_value= -24981;
              imag_value=21194;
            end
    8965  : begin
              real_value= -28766;
              imag_value=15678;
            end
    8966  : begin
              real_value= -31351;
              imag_value=9508;
            end
    8967  : begin
              real_value= -32629;
              imag_value=2942;
            end
    8968  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    8969  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    8970  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    8971  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    8972  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    8973  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    8974  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    8975  : begin
              real_value= -802;
              imag_value=-32750;
            end
    8976  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    8977  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    8978  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    8979  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    8980  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    8981  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    8982  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    8983  : begin
              real_value= 32733;
              imag_value=1338;
            end
    8984  : begin
              real_value= 31779;
              imag_value=7959;
            end
    8985  : begin
              real_value= 29499;
              imag_value=14248;
            end
    8986  : begin
              real_value= 25990;
              imag_value=19943;
            end
    8987  : begin
              real_value= 21399;
              imag_value=24806;
            end
    8988  : begin
              real_value= 15914;
              imag_value=28636;
            end
    8989  : begin
              real_value= 9765;
              imag_value=31271;
            end
    8990  : begin
              real_value= 3210;
              imag_value=32603;
            end
    8991  : begin
              real_value= -3476;
              imag_value=32575;
            end
    8992  : begin
              real_value= -10021;
              imag_value=31191;
            end
    8993  : begin
              real_value= -16148;
              imag_value=28506;
            end
    8994  : begin
              real_value= -21600;
              imag_value=24630;
            end
    8995  : begin
              real_value= -26152;
              imag_value=19729;
            end
    8996  : begin
              real_value= -29615;
              imag_value=14006;
            end
    8997  : begin
              real_value= -31843;
              imag_value=7699;
            end
    8998  : begin
              real_value= -32743;
              imag_value=1070;
            end
    8999  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    9000  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    9001  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    9002  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    9003  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    9004  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    9005  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    9006  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    9007  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    9008  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    9009  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    9010  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    9011  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    9012  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    9013  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    9014  : begin
              real_value= 32603;
              imag_value=3210;
            end
    9015  : begin
              real_value= 31271;
              imag_value=9765;
            end
    9016  : begin
              real_value= 28636;
              imag_value=15914;
            end
    9017  : begin
              real_value= 24806;
              imag_value=21399;
            end
    9018  : begin
              real_value= 19943;
              imag_value=25990;
            end
    9019  : begin
              real_value= 14248;
              imag_value=29499;
            end
    9020  : begin
              real_value= 7959;
              imag_value=31779;
            end
    9021  : begin
              real_value= 1338;
              imag_value=32733;
            end
    9022  : begin
              real_value= -5336;
              imag_value=32323;
            end
    9023  : begin
              real_value= -11790;
              imag_value=30565;
            end
    9024  : begin
              real_value= -17752;
              imag_value=27534;
            end
    9025  : begin
              real_value= -22974;
              imag_value=23354;
            end
    9026  : begin
              real_value= -27240;
              imag_value=18200;
            end
    9027  : begin
              real_value= -30369;
              imag_value=12288;
            end
    9028  : begin
              real_value= -32231;
              imag_value=5864;
            end
    9029  : begin
              real_value= -32750;
              imag_value=-802;
            end
    9030  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    9031  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    9032  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    9033  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    9034  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    9035  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    9036  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    9037  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    9038  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    9039  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    9040  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    9041  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    9042  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    9043  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    9044  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    9045  : begin
              real_value= 32365;
              imag_value=5071;
            end
    9046  : begin
              real_value= 30661;
              imag_value=11539;
            end
    9047  : begin
              real_value= 27678;
              imag_value=17525;
            end
    9048  : begin
              real_value= 23541;
              imag_value=22782;
            end
    9049  : begin
              real_value= 18423;
              imag_value=27090;
            end
    9050  : begin
              real_value= 12537;
              imag_value=30267;
            end
    9051  : begin
              real_value= 6127;
              imag_value=32183;
            end
    9052  : begin
              real_value= -535;
              imag_value=32757;
            end
    9053  : begin
              real_value= -7177;
              imag_value=31965;
            end
    9054  : begin
              real_value= -13520;
              imag_value=29841;
            end
    9055  : begin
              real_value= -19299;
              imag_value=26472;
            end
    9056  : begin
              real_value= -24274;
              imag_value=22001;
            end
    9057  : begin
              real_value= -28236;
              imag_value=16611;
            end
    9058  : begin
              real_value= -31023;
              imag_value=10529;
            end
    9059  : begin
              real_value= -32515;
              imag_value=4009;
            end
    9060  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    9061  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    9062  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    9063  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    9064  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    9065  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    9066  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    9067  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    9068  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    9069  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    9070  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    9071  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    9072  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    9073  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    9074  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    9075  : begin
              real_value= 32759;
              imag_value=267;
            end
    9076  : begin
              real_value= 32022;
              imag_value=6915;
            end
    9077  : begin
              real_value= 29950;
              imag_value=13274;
            end
    9078  : begin
              real_value= 26630;
              imag_value=19081;
            end
    9079  : begin
              real_value= 22199;
              imag_value=24092;
            end
    9080  : begin
              real_value= 16842;
              imag_value=28100;
            end
    9081  : begin
              real_value= 10783;
              imag_value=30935;
            end
    9082  : begin
              real_value= 4275;
              imag_value=32481;
            end
    9083  : begin
              real_value= -2408;
              imag_value=32673;
            end
    9084  : begin
              real_value= -8995;
              imag_value=31501;
            end
    9085  : begin
              real_value= -15206;
              imag_value=29017;
            end
    9086  : begin
              real_value= -20783;
              imag_value=25324;
            end
    9087  : begin
              real_value= -25494;
              imag_value=20575;
            end
    9088  : begin
              real_value= -29142;
              imag_value=14968;
            end
    9089  : begin
              real_value= -31575;
              imag_value=8737;
            end
    9090  : begin
              real_value= -32691;
              imag_value=2142;
            end
    9091  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    9092  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    9093  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    9094  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    9095  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    9096  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    9097  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    9098  : begin
              real_value= 0;
              imag_value=-32760;
            end
    9099  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    9100  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    9101  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    9102  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    9103  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    9104  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    9105  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    9106  : begin
              real_value= 32691;
              imag_value=2142;
            end
    9107  : begin
              real_value= 31575;
              imag_value=8737;
            end
    9108  : begin
              real_value= 29142;
              imag_value=14968;
            end
    9109  : begin
              real_value= 25494;
              imag_value=20575;
            end
    9110  : begin
              real_value= 20783;
              imag_value=25324;
            end
    9111  : begin
              real_value= 15206;
              imag_value=29017;
            end
    9112  : begin
              real_value= 8995;
              imag_value=31501;
            end
    9113  : begin
              real_value= 2408;
              imag_value=32673;
            end
    9114  : begin
              real_value= -4275;
              imag_value=32481;
            end
    9115  : begin
              real_value= -10783;
              imag_value=30935;
            end
    9116  : begin
              real_value= -16842;
              imag_value=28100;
            end
    9117  : begin
              real_value= -22199;
              imag_value=24092;
            end
    9118  : begin
              real_value= -26630;
              imag_value=19081;
            end
    9119  : begin
              real_value= -29950;
              imag_value=13274;
            end
    9120  : begin
              real_value= -32022;
              imag_value=6915;
            end
    9121  : begin
              real_value= -32759;
              imag_value=267;
            end
    9122  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    9123  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    9124  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    9125  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    9126  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    9127  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    9128  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    9129  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    9130  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    9131  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    9132  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    9133  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    9134  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    9135  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    9136  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    9137  : begin
              real_value= 32515;
              imag_value=4009;
            end
    9138  : begin
              real_value= 31023;
              imag_value=10529;
            end
    9139  : begin
              real_value= 28236;
              imag_value=16611;
            end
    9140  : begin
              real_value= 24274;
              imag_value=22001;
            end
    9141  : begin
              real_value= 19299;
              imag_value=26472;
            end
    9142  : begin
              real_value= 13520;
              imag_value=29841;
            end
    9143  : begin
              real_value= 7177;
              imag_value=31965;
            end
    9144  : begin
              real_value= 535;
              imag_value=32757;
            end
    9145  : begin
              real_value= -6127;
              imag_value=32183;
            end
    9146  : begin
              real_value= -12537;
              imag_value=30267;
            end
    9147  : begin
              real_value= -18423;
              imag_value=27090;
            end
    9148  : begin
              real_value= -23541;
              imag_value=22782;
            end
    9149  : begin
              real_value= -27678;
              imag_value=17525;
            end
    9150  : begin
              real_value= -30661;
              imag_value=11539;
            end
    9151  : begin
              real_value= -32365;
              imag_value=5071;
            end
    9152  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    9153  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    9154  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    9155  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    9156  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    9157  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    9158  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    9159  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    9160  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    9161  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    9162  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    9163  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    9164  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    9165  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    9166  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    9167  : begin
              real_value= 32750;
              imag_value=-802;
            end
    9168  : begin
              real_value= 32231;
              imag_value=5864;
            end
    9169  : begin
              real_value= 30369;
              imag_value=12288;
            end
    9170  : begin
              real_value= 27240;
              imag_value=18200;
            end
    9171  : begin
              real_value= 22974;
              imag_value=23354;
            end
    9172  : begin
              real_value= 17752;
              imag_value=27534;
            end
    9173  : begin
              real_value= 11790;
              imag_value=30565;
            end
    9174  : begin
              real_value= 5336;
              imag_value=32323;
            end
    9175  : begin
              real_value= -1338;
              imag_value=32733;
            end
    9176  : begin
              real_value= -7959;
              imag_value=31779;
            end
    9177  : begin
              real_value= -14248;
              imag_value=29499;
            end
    9178  : begin
              real_value= -19943;
              imag_value=25990;
            end
    9179  : begin
              real_value= -24806;
              imag_value=21399;
            end
    9180  : begin
              real_value= -28636;
              imag_value=15914;
            end
    9181  : begin
              real_value= -31271;
              imag_value=9765;
            end
    9182  : begin
              real_value= -32603;
              imag_value=3210;
            end
    9183  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    9184  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    9185  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    9186  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    9187  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    9188  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    9189  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    9190  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    9191  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    9192  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    9193  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    9194  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    9195  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    9196  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    9197  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    9198  : begin
              real_value= 32743;
              imag_value=1070;
            end
    9199  : begin
              real_value= 31843;
              imag_value=7699;
            end
    9200  : begin
              real_value= 29615;
              imag_value=14006;
            end
    9201  : begin
              real_value= 26152;
              imag_value=19729;
            end
    9202  : begin
              real_value= 21600;
              imag_value=24630;
            end
    9203  : begin
              real_value= 16148;
              imag_value=28506;
            end
    9204  : begin
              real_value= 10021;
              imag_value=31191;
            end
    9205  : begin
              real_value= 3476;
              imag_value=32575;
            end
    9206  : begin
              real_value= -3210;
              imag_value=32603;
            end
    9207  : begin
              real_value= -9765;
              imag_value=31271;
            end
    9208  : begin
              real_value= -15914;
              imag_value=28636;
            end
    9209  : begin
              real_value= -21399;
              imag_value=24806;
            end
    9210  : begin
              real_value= -25990;
              imag_value=19943;
            end
    9211  : begin
              real_value= -29499;
              imag_value=14248;
            end
    9212  : begin
              real_value= -31779;
              imag_value=7959;
            end
    9213  : begin
              real_value= -32733;
              imag_value=1338;
            end
    9214  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    9215  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    9216  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    9217  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    9218  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    9219  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    9220  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    9221  : begin
              real_value= 802;
              imag_value=-32750;
            end
    9222  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    9223  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    9224  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    9225  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    9226  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    9227  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    9228  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    9229  : begin
              real_value= 32629;
              imag_value=2942;
            end
    9230  : begin
              real_value= 31351;
              imag_value=9508;
            end
    9231  : begin
              real_value= 28766;
              imag_value=15678;
            end
    9232  : begin
              real_value= 24981;
              imag_value=21194;
            end
    9233  : begin
              real_value= 20154;
              imag_value=25826;
            end
    9234  : begin
              real_value= 14489;
              imag_value=29382;
            end
    9235  : begin
              real_value= 8219;
              imag_value=31713;
            end
    9236  : begin
              real_value= 1606;
              imag_value=32721;
            end
    9237  : begin
              real_value= -5071;
              imag_value=32365;
            end
    9238  : begin
              real_value= -11539;
              imag_value=30661;
            end
    9239  : begin
              real_value= -17525;
              imag_value=27678;
            end
    9240  : begin
              real_value= -22782;
              imag_value=23541;
            end
    9241  : begin
              real_value= -27090;
              imag_value=18423;
            end
    9242  : begin
              real_value= -30267;
              imag_value=12537;
            end
    9243  : begin
              real_value= -32183;
              imag_value=6127;
            end
    9244  : begin
              real_value= -32757;
              imag_value=-535;
            end
    9245  : begin
              real_value= -31965;
              imag_value=-7177;
            end
    9246  : begin
              real_value= -29841;
              imag_value=-13520;
            end
    9247  : begin
              real_value= -26472;
              imag_value=-19299;
            end
    9248  : begin
              real_value= -22001;
              imag_value=-24274;
            end
    9249  : begin
              real_value= -16611;
              imag_value=-28236;
            end
    9250  : begin
              real_value= -10529;
              imag_value=-31023;
            end
    9251  : begin
              real_value= -4009;
              imag_value=-32515;
            end
    9252  : begin
              real_value= 2676;
              imag_value=-32651;
            end
    9253  : begin
              real_value= 9253;
              imag_value=-31426;
            end
    9254  : begin
              real_value= 15442;
              imag_value=-28892;
            end
    9255  : begin
              real_value= 20988;
              imag_value=-25154;
            end
    9256  : begin
              real_value= 25661;
              imag_value=-20365;
            end
    9257  : begin
              real_value= 29263;
              imag_value=-14728;
            end
    9258  : begin
              real_value= 31645;
              imag_value=-8477;
            end
    9259  : begin
              real_value= 32707;
              imag_value=-1874;
            end
    9260  : begin
              real_value= 32407;
              imag_value=4806;
            end
    9261  : begin
              real_value= 30755;
              imag_value=11289;
            end
    9262  : begin
              real_value= 27820;
              imag_value=17299;
            end
    9263  : begin
              real_value= 23726;
              imag_value=22589;
            end
    9264  : begin
              real_value= 18644;
              imag_value=26938;
            end
    9265  : begin
              real_value= 12784;
              imag_value=30163;
            end
    9266  : begin
              real_value= 6390;
              imag_value=32131;
            end
    9267  : begin
              real_value= -267;
              imag_value=32759;
            end
    9268  : begin
              real_value= -6915;
              imag_value=32022;
            end
    9269  : begin
              real_value= -13274;
              imag_value=29950;
            end
    9270  : begin
              real_value= -19081;
              imag_value=26630;
            end
    9271  : begin
              real_value= -24092;
              imag_value=22199;
            end
    9272  : begin
              real_value= -28100;
              imag_value=16842;
            end
    9273  : begin
              real_value= -30935;
              imag_value=10783;
            end
    9274  : begin
              real_value= -32481;
              imag_value=4275;
            end
    9275  : begin
              real_value= -32673;
              imag_value=-2408;
            end
    9276  : begin
              real_value= -31501;
              imag_value=-8995;
            end
    9277  : begin
              real_value= -29017;
              imag_value=-15206;
            end
    9278  : begin
              real_value= -25324;
              imag_value=-20783;
            end
    9279  : begin
              real_value= -20575;
              imag_value=-25494;
            end
    9280  : begin
              real_value= -14968;
              imag_value=-29142;
            end
    9281  : begin
              real_value= -8737;
              imag_value=-31575;
            end
    9282  : begin
              real_value= -2142;
              imag_value=-32691;
            end
    9283  : begin
              real_value= 4540;
              imag_value=-32445;
            end
    9284  : begin
              real_value= 11036;
              imag_value=-30846;
            end
    9285  : begin
              real_value= 17072;
              imag_value=-27961;
            end
    9286  : begin
              real_value= 22395;
              imag_value=-23911;
            end
    9287  : begin
              real_value= 26784;
              imag_value=-18863;
            end
    9288  : begin
              real_value= 30057;
              imag_value=-13030;
            end
    9289  : begin
              real_value= 32077;
              imag_value=-6654;
            end
    9290  : begin
              real_value= 32760;
              imag_value=0;
            end
    9291  : begin
              real_value= 32077;
              imag_value=6654;
            end
    9292  : begin
              real_value= 30057;
              imag_value=13030;
            end
    9293  : begin
              real_value= 26784;
              imag_value=18863;
            end
    9294  : begin
              real_value= 22395;
              imag_value=23911;
            end
    9295  : begin
              real_value= 17072;
              imag_value=27961;
            end
    9296  : begin
              real_value= 11036;
              imag_value=30846;
            end
    9297  : begin
              real_value= 4540;
              imag_value=32445;
            end
    9298  : begin
              real_value= -2142;
              imag_value=32691;
            end
    9299  : begin
              real_value= -8737;
              imag_value=31575;
            end
    9300  : begin
              real_value= -14968;
              imag_value=29142;
            end
    9301  : begin
              real_value= -20575;
              imag_value=25494;
            end
    9302  : begin
              real_value= -25324;
              imag_value=20783;
            end
    9303  : begin
              real_value= -29017;
              imag_value=15206;
            end
    9304  : begin
              real_value= -31501;
              imag_value=8995;
            end
    9305  : begin
              real_value= -32673;
              imag_value=2408;
            end
    9306  : begin
              real_value= -32481;
              imag_value=-4275;
            end
    9307  : begin
              real_value= -30935;
              imag_value=-10783;
            end
    9308  : begin
              real_value= -28100;
              imag_value=-16842;
            end
    9309  : begin
              real_value= -24092;
              imag_value=-22199;
            end
    9310  : begin
              real_value= -19081;
              imag_value=-26630;
            end
    9311  : begin
              real_value= -13274;
              imag_value=-29950;
            end
    9312  : begin
              real_value= -6915;
              imag_value=-32022;
            end
    9313  : begin
              real_value= -267;
              imag_value=-32759;
            end
    9314  : begin
              real_value= 6390;
              imag_value=-32131;
            end
    9315  : begin
              real_value= 12784;
              imag_value=-30163;
            end
    9316  : begin
              real_value= 18644;
              imag_value=-26938;
            end
    9317  : begin
              real_value= 23726;
              imag_value=-22589;
            end
    9318  : begin
              real_value= 27820;
              imag_value=-17299;
            end
    9319  : begin
              real_value= 30755;
              imag_value=-11289;
            end
    9320  : begin
              real_value= 32407;
              imag_value=-4806;
            end
    9321  : begin
              real_value= 32707;
              imag_value=1874;
            end
    9322  : begin
              real_value= 31645;
              imag_value=8477;
            end
    9323  : begin
              real_value= 29263;
              imag_value=14728;
            end
    9324  : begin
              real_value= 25661;
              imag_value=20365;
            end
    9325  : begin
              real_value= 20988;
              imag_value=25154;
            end
    9326  : begin
              real_value= 15442;
              imag_value=28892;
            end
    9327  : begin
              real_value= 9253;
              imag_value=31426;
            end
    9328  : begin
              real_value= 2676;
              imag_value=32651;
            end
    9329  : begin
              real_value= -4009;
              imag_value=32515;
            end
    9330  : begin
              real_value= -10529;
              imag_value=31023;
            end
    9331  : begin
              real_value= -16611;
              imag_value=28236;
            end
    9332  : begin
              real_value= -22001;
              imag_value=24274;
            end
    9333  : begin
              real_value= -26472;
              imag_value=19299;
            end
    9334  : begin
              real_value= -29841;
              imag_value=13520;
            end
    9335  : begin
              real_value= -31965;
              imag_value=7177;
            end
    9336  : begin
              real_value= -32757;
              imag_value=535;
            end
    9337  : begin
              real_value= -32183;
              imag_value=-6127;
            end
    9338  : begin
              real_value= -30267;
              imag_value=-12537;
            end
    9339  : begin
              real_value= -27090;
              imag_value=-18423;
            end
    9340  : begin
              real_value= -22782;
              imag_value=-23541;
            end
    9341  : begin
              real_value= -17525;
              imag_value=-27678;
            end
    9342  : begin
              real_value= -11539;
              imag_value=-30661;
            end
    9343  : begin
              real_value= -5071;
              imag_value=-32365;
            end
    9344  : begin
              real_value= 1606;
              imag_value=-32721;
            end
    9345  : begin
              real_value= 8219;
              imag_value=-31713;
            end
    9346  : begin
              real_value= 14489;
              imag_value=-29382;
            end
    9347  : begin
              real_value= 20154;
              imag_value=-25826;
            end
    9348  : begin
              real_value= 24981;
              imag_value=-21194;
            end
    9349  : begin
              real_value= 28766;
              imag_value=-15678;
            end
    9350  : begin
              real_value= 31351;
              imag_value=-9508;
            end
    9351  : begin
              real_value= 32629;
              imag_value=-2942;
            end
    9352  : begin
              real_value= 32547;
              imag_value=3742;
            end
    9353  : begin
              real_value= 31107;
              imag_value=10275;
            end
    9354  : begin
              real_value= 28371;
              imag_value=16380;
            end
    9355  : begin
              real_value= 24453;
              imag_value=21801;
            end
    9356  : begin
              real_value= 19515;
              imag_value=26314;
            end
    9357  : begin
              real_value= 13764;
              imag_value=29729;
            end
    9358  : begin
              real_value= 7438;
              imag_value=31905;
            end
    9359  : begin
              real_value= 802;
              imag_value=32750;
            end
    9360  : begin
              real_value= -5864;
              imag_value=32231;
            end
    9361  : begin
              real_value= -12288;
              imag_value=30369;
            end
    9362  : begin
              real_value= -18200;
              imag_value=27240;
            end
    9363  : begin
              real_value= -23354;
              imag_value=22974;
            end
    9364  : begin
              real_value= -27534;
              imag_value=17752;
            end
    9365  : begin
              real_value= -30565;
              imag_value=11790;
            end
    9366  : begin
              real_value= -32323;
              imag_value=5336;
            end
    9367  : begin
              real_value= -32733;
              imag_value=-1338;
            end
    9368  : begin
              real_value= -31779;
              imag_value=-7959;
            end
    9369  : begin
              real_value= -29499;
              imag_value=-14248;
            end
    9370  : begin
              real_value= -25990;
              imag_value=-19943;
            end
    9371  : begin
              real_value= -21399;
              imag_value=-24806;
            end
    9372  : begin
              real_value= -15914;
              imag_value=-28636;
            end
    9373  : begin
              real_value= -9765;
              imag_value=-31271;
            end
    9374  : begin
              real_value= -3210;
              imag_value=-32603;
            end
    9375  : begin
              real_value= 3476;
              imag_value=-32575;
            end
    9376  : begin
              real_value= 10021;
              imag_value=-31191;
            end
    9377  : begin
              real_value= 16148;
              imag_value=-28506;
            end
    9378  : begin
              real_value= 21600;
              imag_value=-24630;
            end
    9379  : begin
              real_value= 26152;
              imag_value=-19729;
            end
    9380  : begin
              real_value= 29615;
              imag_value=-14006;
            end
    9381  : begin
              real_value= 31843;
              imag_value=-7699;
            end
    9382  : begin
              real_value= 32743;
              imag_value=-1070;
            end
    9383  : begin
              real_value= 32278;
              imag_value=5599;
            end
    9384  : begin
              real_value= 30468;
              imag_value=12039;
            end
    9385  : begin
              real_value= 27387;
              imag_value=17977;
            end
    9386  : begin
              real_value= 23165;
              imag_value=23165;
            end
    9387  : begin
              real_value= 17977;
              imag_value=27387;
            end
    9388  : begin
              real_value= 12039;
              imag_value=30468;
            end
    9389  : begin
              real_value= 5599;
              imag_value=32278;
            end
    9390  : begin
              real_value= -1070;
              imag_value=32743;
            end
    9391  : begin
              real_value= -7699;
              imag_value=31843;
            end
    9392  : begin
              real_value= -14006;
              imag_value=29615;
            end
    9393  : begin
              real_value= -19729;
              imag_value=26152;
            end
    9394  : begin
              real_value= -24630;
              imag_value=21600;
            end
    9395  : begin
              real_value= -28506;
              imag_value=16148;
            end
    9396  : begin
              real_value= -31191;
              imag_value=10021;
            end
    9397  : begin
              real_value= -32575;
              imag_value=3476;
            end
    9398  : begin
              real_value= -32603;
              imag_value=-3210;
            end
    9399  : begin
              real_value= -31271;
              imag_value=-9765;
            end
    9400  : begin
              real_value= -28636;
              imag_value=-15914;
            end
    9401  : begin
              real_value= -24806;
              imag_value=-21399;
            end
    9402  : begin
              real_value= -19943;
              imag_value=-25990;
            end
    9403  : begin
              real_value= -14248;
              imag_value=-29499;
            end
    9404  : begin
              real_value= -7959;
              imag_value=-31779;
            end
    9405  : begin
              real_value= -1338;
              imag_value=-32733;
            end
    9406  : begin
              real_value= 5336;
              imag_value=-32323;
            end
    9407  : begin
              real_value= 11790;
              imag_value=-30565;
            end
    9408  : begin
              real_value= 17752;
              imag_value=-27534;
            end
    9409  : begin
              real_value= 22974;
              imag_value=-23354;
            end
    9410  : begin
              real_value= 27240;
              imag_value=-18200;
            end
    9411  : begin
              real_value= 30369;
              imag_value=-12288;
            end
    9412  : begin
              real_value= 32231;
              imag_value=-5864;
            end
    9413  : begin
              real_value= 32750;
              imag_value=802;
            end
    9414  : begin
              real_value= 31905;
              imag_value=7438;
            end
    9415  : begin
              real_value= 29729;
              imag_value=13764;
            end
    9416  : begin
              real_value= 26314;
              imag_value=19515;
            end
    9417  : begin
              real_value= 21801;
              imag_value=24453;
            end
    9418  : begin
              real_value= 16380;
              imag_value=28371;
            end
    9419  : begin
              real_value= 10275;
              imag_value=31107;
            end
    9420  : begin
              real_value= 3742;
              imag_value=32547;
            end
    9421  : begin
              real_value= -2942;
              imag_value=32629;
            end
    9422  : begin
              real_value= -9508;
              imag_value=31351;
            end
    9423  : begin
              real_value= -15678;
              imag_value=28766;
            end
    9424  : begin
              real_value= -21194;
              imag_value=24981;
            end
    9425  : begin
              real_value= -25826;
              imag_value=20154;
            end
    9426  : begin
              real_value= -29382;
              imag_value=14489;
            end
    9427  : begin
              real_value= -31713;
              imag_value=8219;
            end
    9428  : begin
              real_value= -32721;
              imag_value=1606;
            end
    9429  : begin
              real_value= -32365;
              imag_value=-5071;
            end
    9430  : begin
              real_value= -30661;
              imag_value=-11539;
            end
    9431  : begin
              real_value= -27678;
              imag_value=-17525;
            end
    9432  : begin
              real_value= -23541;
              imag_value=-22782;
            end
    9433  : begin
              real_value= -18423;
              imag_value=-27090;
            end
    9434  : begin
              real_value= -12537;
              imag_value=-30267;
            end
    9435  : begin
              real_value= -6127;
              imag_value=-32183;
            end
    9436  : begin
              real_value= 535;
              imag_value=-32757;
            end
    9437  : begin
              real_value= 7177;
              imag_value=-31965;
            end
    9438  : begin
              real_value= 13520;
              imag_value=-29841;
            end
    9439  : begin
              real_value= 19299;
              imag_value=-26472;
            end
    9440  : begin
              real_value= 24274;
              imag_value=-22001;
            end
    9441  : begin
              real_value= 28236;
              imag_value=-16611;
            end
    9442  : begin
              real_value= 31023;
              imag_value=-10529;
            end
    9443  : begin
              real_value= 32515;
              imag_value=-4009;
            end
    9444  : begin
              real_value= 32651;
              imag_value=2676;
            end
    9445  : begin
              real_value= 31426;
              imag_value=9253;
            end
    9446  : begin
              real_value= 28892;
              imag_value=15442;
            end
    9447  : begin
              real_value= 25154;
              imag_value=20988;
            end
    9448  : begin
              real_value= 20365;
              imag_value=25661;
            end
    9449  : begin
              real_value= 14728;
              imag_value=29263;
            end
    9450  : begin
              real_value= 8477;
              imag_value=31645;
            end
    9451  : begin
              real_value= 1874;
              imag_value=32707;
            end
    9452  : begin
              real_value= -4806;
              imag_value=32407;
            end
    9453  : begin
              real_value= -11289;
              imag_value=30755;
            end
    9454  : begin
              real_value= -17299;
              imag_value=27820;
            end
    9455  : begin
              real_value= -22589;
              imag_value=23726;
            end
    9456  : begin
              real_value= -26938;
              imag_value=18644;
            end
    9457  : begin
              real_value= -30163;
              imag_value=12784;
            end
    9458  : begin
              real_value= -32131;
              imag_value=6390;
            end
    9459  : begin
              real_value= -32759;
              imag_value=-267;
            end
    9460  : begin
              real_value= -32022;
              imag_value=-6915;
            end
    9461  : begin
              real_value= -29950;
              imag_value=-13274;
            end
    9462  : begin
              real_value= -26630;
              imag_value=-19081;
            end
    9463  : begin
              real_value= -22199;
              imag_value=-24092;
            end
    9464  : begin
              real_value= -16842;
              imag_value=-28100;
            end
    9465  : begin
              real_value= -10783;
              imag_value=-30935;
            end
    9466  : begin
              real_value= -4275;
              imag_value=-32481;
            end
    9467  : begin
              real_value= 2408;
              imag_value=-32673;
            end
    9468  : begin
              real_value= 8995;
              imag_value=-31501;
            end
    9469  : begin
              real_value= 15206;
              imag_value=-29017;
            end
    9470  : begin
              real_value= 20783;
              imag_value=-25324;
            end
    9471  : begin
              real_value= 25494;
              imag_value=-20575;
            end
    9472  : begin
              real_value= 29142;
              imag_value=-14968;
            end
    9473  : begin
              real_value= 31575;
              imag_value=-8737;
            end
    9474  : begin
              real_value= 32691;
              imag_value=-2142;
            end
    9475  : begin
              real_value= 32445;
              imag_value=4540;
            end
    9476  : begin
              real_value= 30846;
              imag_value=11036;
            end
    9477  : begin
              real_value= 27961;
              imag_value=17072;
            end
    9478  : begin
              real_value= 23911;
              imag_value=22395;
            end
    9479  : begin
              real_value= 18863;
              imag_value=26784;
            end
    9480  : begin
              real_value= 13030;
              imag_value=30057;
            end
    9481  : begin
              real_value= 6654;
              imag_value=32077;
            end
    9482  : begin
              real_value= 0;
              imag_value=32760;
            end
    9483  : begin
              real_value= -6654;
              imag_value=32077;
            end
    9484  : begin
              real_value= -13030;
              imag_value=30057;
            end
    9485  : begin
              real_value= -18863;
              imag_value=26784;
            end
    9486  : begin
              real_value= -23911;
              imag_value=22395;
            end
    9487  : begin
              real_value= -27961;
              imag_value=17072;
            end
    9488  : begin
              real_value= -30846;
              imag_value=11036;
            end
    9489  : begin
              real_value= -32445;
              imag_value=4540;
            end
    9490  : begin
              real_value= -32691;
              imag_value=-2142;
            end
    9491  : begin
              real_value= -31575;
              imag_value=-8737;
            end
    9492  : begin
              real_value= -29142;
              imag_value=-14968;
            end
    9493  : begin
              real_value= -25494;
              imag_value=-20575;
            end
    9494  : begin
              real_value= -20783;
              imag_value=-25324;
            end
    9495  : begin
              real_value= -15206;
              imag_value=-29017;
            end
    9496  : begin
              real_value= -8995;
              imag_value=-31501;
            end
    9497  : begin
              real_value= -2408;
              imag_value=-32673;
            end
    9498  : begin
              real_value= 4275;
              imag_value=-32481;
            end
    9499  : begin
              real_value= 10783;
              imag_value=-30935;
            end
    9500  : begin
              real_value= 16842;
              imag_value=-28100;
            end
    9501  : begin
              real_value= 22199;
              imag_value=-24092;
            end
    9502  : begin
              real_value= 26630;
              imag_value=-19081;
            end
    9503  : begin
              real_value= 29950;
              imag_value=-13274;
            end
    9504  : begin
              real_value= 32022;
              imag_value=-6915;
            end
    9505  : begin
              real_value= 32759;
              imag_value=-267;
            end
    9506  : begin
              real_value= 32131;
              imag_value=6390;
            end
    9507  : begin
              real_value= 30163;
              imag_value=12784;
            end
    9508  : begin
              real_value= 26938;
              imag_value=18644;
            end
    9509  : begin
              real_value= 22589;
              imag_value=23726;
            end
    9510  : begin
              real_value= 17299;
              imag_value=27820;
            end
    9511  : begin
              real_value= 11289;
              imag_value=30755;
            end
    9512  : begin
              real_value= 4806;
              imag_value=32407;
            end
    9513  : begin
              real_value= -1874;
              imag_value=32707;
            end
    9514  : begin
              real_value= -8477;
              imag_value=31645;
            end
    9515  : begin
              real_value= -14728;
              imag_value=29263;
            end
    9516  : begin
              real_value= -20365;
              imag_value=25661;
            end
    9517  : begin
              real_value= -25154;
              imag_value=20988;
            end
    9518  : begin
              real_value= -28892;
              imag_value=15442;
            end
    9519  : begin
              real_value= -31426;
              imag_value=9253;
            end
    9520  : begin
              real_value= -32651;
              imag_value=2676;
            end
    9521  : begin
              real_value= -32515;
              imag_value=-4009;
            end
    9522  : begin
              real_value= -31023;
              imag_value=-10529;
            end
    9523  : begin
              real_value= -28236;
              imag_value=-16611;
            end
    9524  : begin
              real_value= -24274;
              imag_value=-22001;
            end
    9525  : begin
              real_value= -19299;
              imag_value=-26472;
            end
    9526  : begin
              real_value= -13520;
              imag_value=-29841;
            end
    9527  : begin
              real_value= -7177;
              imag_value=-31965;
            end
    9528  : begin
              real_value= -535;
              imag_value=-32757;
            end
    9529  : begin
              real_value= 6127;
              imag_value=-32183;
            end
    9530  : begin
              real_value= 12537;
              imag_value=-30267;
            end
    9531  : begin
              real_value= 18423;
              imag_value=-27090;
            end
    9532  : begin
              real_value= 23541;
              imag_value=-22782;
            end
    9533  : begin
              real_value= 27678;
              imag_value=-17525;
            end
    9534  : begin
              real_value= 30661;
              imag_value=-11539;
            end
    9535  : begin
              real_value= 32365;
              imag_value=-5071;
            end
    9536  : begin
              real_value= 32721;
              imag_value=1606;
            end
    9537  : begin
              real_value= 31713;
              imag_value=8219;
            end
    9538  : begin
              real_value= 29382;
              imag_value=14489;
            end
    9539  : begin
              real_value= 25826;
              imag_value=20154;
            end
    9540  : begin
              real_value= 21194;
              imag_value=24981;
            end
    9541  : begin
              real_value= 15678;
              imag_value=28766;
            end
    9542  : begin
              real_value= 9508;
              imag_value=31351;
            end
    9543  : begin
              real_value= 2942;
              imag_value=32629;
            end
    9544  : begin
              real_value= -3742;
              imag_value=32547;
            end
    9545  : begin
              real_value= -10275;
              imag_value=31107;
            end
    9546  : begin
              real_value= -16380;
              imag_value=28371;
            end
    9547  : begin
              real_value= -21801;
              imag_value=24453;
            end
    9548  : begin
              real_value= -26314;
              imag_value=19515;
            end
    9549  : begin
              real_value= -29729;
              imag_value=13764;
            end
    9550  : begin
              real_value= -31905;
              imag_value=7438;
            end
    9551  : begin
              real_value= -32750;
              imag_value=802;
            end
    9552  : begin
              real_value= -32231;
              imag_value=-5864;
            end
    9553  : begin
              real_value= -30369;
              imag_value=-12288;
            end
    9554  : begin
              real_value= -27240;
              imag_value=-18200;
            end
    9555  : begin
              real_value= -22974;
              imag_value=-23354;
            end
    9556  : begin
              real_value= -17752;
              imag_value=-27534;
            end
    9557  : begin
              real_value= -11790;
              imag_value=-30565;
            end
    9558  : begin
              real_value= -5336;
              imag_value=-32323;
            end
    9559  : begin
              real_value= 1338;
              imag_value=-32733;
            end
    9560  : begin
              real_value= 7959;
              imag_value=-31779;
            end
    9561  : begin
              real_value= 14248;
              imag_value=-29499;
            end
    9562  : begin
              real_value= 19943;
              imag_value=-25990;
            end
    9563  : begin
              real_value= 24806;
              imag_value=-21399;
            end
    9564  : begin
              real_value= 28636;
              imag_value=-15914;
            end
    9565  : begin
              real_value= 31271;
              imag_value=-9765;
            end
    9566  : begin
              real_value= 32603;
              imag_value=-3210;
            end
    9567  : begin
              real_value= 32575;
              imag_value=3476;
            end
    9568  : begin
              real_value= 31191;
              imag_value=10021;
            end
    9569  : begin
              real_value= 28506;
              imag_value=16148;
            end
    9570  : begin
              real_value= 24630;
              imag_value=21600;
            end
    9571  : begin
              real_value= 19729;
              imag_value=26152;
            end
    9572  : begin
              real_value= 14006;
              imag_value=29615;
            end
    9573  : begin
              real_value= 7699;
              imag_value=31843;
            end
    9574  : begin
              real_value= 1070;
              imag_value=32743;
            end
    9575  : begin
              real_value= -5599;
              imag_value=32278;
            end
    9576  : begin
              real_value= -12039;
              imag_value=30468;
            end
    9577  : begin
              real_value= -17977;
              imag_value=27387;
            end
    9578  : begin
              real_value= -23165;
              imag_value=23165;
            end
    9579  : begin
              real_value= -27387;
              imag_value=17977;
            end
    9580  : begin
              real_value= -30468;
              imag_value=12039;
            end
    9581  : begin
              real_value= -32278;
              imag_value=5599;
            end
    9582  : begin
              real_value= -32743;
              imag_value=-1070;
            end
    9583  : begin
              real_value= -31843;
              imag_value=-7699;
            end
    9584  : begin
              real_value= -29615;
              imag_value=-14006;
            end
    9585  : begin
              real_value= -26152;
              imag_value=-19729;
            end
    9586  : begin
              real_value= -21600;
              imag_value=-24630;
            end
    9587  : begin
              real_value= -16148;
              imag_value=-28506;
            end
    9588  : begin
              real_value= -10021;
              imag_value=-31191;
            end
    9589  : begin
              real_value= -3476;
              imag_value=-32575;
            end
    9590  : begin
              real_value= 3210;
              imag_value=-32603;
            end
    9591  : begin
              real_value= 9765;
              imag_value=-31271;
            end
    9592  : begin
              real_value= 15914;
              imag_value=-28636;
            end
    9593  : begin
              real_value= 21399;
              imag_value=-24806;
            end
    9594  : begin
              real_value= 25990;
              imag_value=-19943;
            end
    9595  : begin
              real_value= 29499;
              imag_value=-14248;
            end
    9596  : begin
              real_value= 31779;
              imag_value=-7959;
            end
    9597  : begin
              real_value= 32733;
              imag_value=-1338;
            end
    9598  : begin
              real_value= 32323;
              imag_value=5336;
            end
    9599  : begin
              real_value= 30565;
              imag_value=11790;
            end
    9600  : begin
              real_value= 27534;
              imag_value=17752;
            end
    9601  : begin
              real_value= 23354;
              imag_value=22974;
            end
    9602  : begin
              real_value= 18200;
              imag_value=27240;
            end
    9603  : begin
              real_value= 12288;
              imag_value=30369;
            end
    9604  : begin
              real_value= 5864;
              imag_value=32231;
            end
    9605  : begin
              real_value= -802;
              imag_value=32750;
            end
    9606  : begin
              real_value= -7438;
              imag_value=31905;
            end
    9607  : begin
              real_value= -13764;
              imag_value=29729;
            end
    9608  : begin
              real_value= -19515;
              imag_value=26314;
            end
    9609  : begin
              real_value= -24453;
              imag_value=21801;
            end
    9610  : begin
              real_value= -28371;
              imag_value=16380;
            end
    9611  : begin
              real_value= -31107;
              imag_value=10275;
            end
    9612  : begin
              real_value= -32547;
              imag_value=3742;
            end
    9613  : begin
              real_value= -32629;
              imag_value=-2942;
            end
    9614  : begin
              real_value= -31351;
              imag_value=-9508;
            end
    9615  : begin
              real_value= -28766;
              imag_value=-15678;
            end
    9616  : begin
              real_value= -24981;
              imag_value=-21194;
            end
    9617  : begin
              real_value= -20154;
              imag_value=-25826;
            end
    9618  : begin
              real_value= -14489;
              imag_value=-29382;
            end
    9619  : begin
              real_value= -8219;
              imag_value=-31713;
            end
    9620  : begin
              real_value= -1606;
              imag_value=-32721;
            end
    9621  : begin
              real_value= 5071;
              imag_value=-32365;
            end
    9622  : begin
              real_value= 11539;
              imag_value=-30661;
            end
    9623  : begin
              real_value= 17525;
              imag_value=-27678;
            end
    9624  : begin
              real_value= 22782;
              imag_value=-23541;
            end
    9625  : begin
              real_value= 27090;
              imag_value=-18423;
            end
    9626  : begin
              real_value= 30267;
              imag_value=-12537;
            end
    9627  : begin
              real_value= 32183;
              imag_value=-6127;
            end
    9628  : begin
              real_value= 32757;
              imag_value=535;
            end
    9629  : begin
              real_value= 31965;
              imag_value=7177;
            end
    9630  : begin
              real_value= 29841;
              imag_value=13520;
            end
    9631  : begin
              real_value= 26472;
              imag_value=19299;
            end
    9632  : begin
              real_value= 22001;
              imag_value=24274;
            end
    9633  : begin
              real_value= 16611;
              imag_value=28236;
            end
    9634  : begin
              real_value= 10529;
              imag_value=31023;
            end
    9635  : begin
              real_value= 4009;
              imag_value=32515;
            end
    9636  : begin
              real_value= -2676;
              imag_value=32651;
            end
    9637  : begin
              real_value= -9253;
              imag_value=31426;
            end
    9638  : begin
              real_value= -15442;
              imag_value=28892;
            end
    9639  : begin
              real_value= -20988;
              imag_value=25154;
            end
    9640  : begin
              real_value= -25661;
              imag_value=20365;
            end
    9641  : begin
              real_value= -29263;
              imag_value=14728;
            end
    9642  : begin
              real_value= -31645;
              imag_value=8477;
            end
    9643  : begin
              real_value= -32707;
              imag_value=1874;
            end
    9644  : begin
              real_value= -32407;
              imag_value=-4806;
            end
    9645  : begin
              real_value= -30755;
              imag_value=-11289;
            end
    9646  : begin
              real_value= -27820;
              imag_value=-17299;
            end
    9647  : begin
              real_value= -23726;
              imag_value=-22589;
            end
    9648  : begin
              real_value= -18644;
              imag_value=-26938;
            end
    9649  : begin
              real_value= -12784;
              imag_value=-30163;
            end
    9650  : begin
              real_value= -6390;
              imag_value=-32131;
            end
    9651  : begin
              real_value= 267;
              imag_value=-32759;
            end
    9652  : begin
              real_value= 6915;
              imag_value=-32022;
            end
    9653  : begin
              real_value= 13274;
              imag_value=-29950;
            end
    9654  : begin
              real_value= 19081;
              imag_value=-26630;
            end
    9655  : begin
              real_value= 24092;
              imag_value=-22199;
            end
    9656  : begin
              real_value= 28100;
              imag_value=-16842;
            end
    9657  : begin
              real_value= 30935;
              imag_value=-10783;
            end
    9658  : begin
              real_value= 32481;
              imag_value=-4275;
            end
    9659  : begin
              real_value= 32673;
              imag_value=2408;
            end
    9660  : begin
              real_value= 31501;
              imag_value=8995;
            end
    9661  : begin
              real_value= 29017;
              imag_value=15206;
            end
    9662  : begin
              real_value= 25324;
              imag_value=20783;
            end
    9663  : begin
              real_value= 20575;
              imag_value=25494;
            end
    9664  : begin
              real_value= 14968;
              imag_value=29142;
            end
    9665  : begin
              real_value= 8737;
              imag_value=31575;
            end
    9666  : begin
              real_value= 2142;
              imag_value=32691;
            end
    9667  : begin
              real_value= -4540;
              imag_value=32445;
            end
    9668  : begin
              real_value= -11036;
              imag_value=30846;
            end
    9669  : begin
              real_value= -17072;
              imag_value=27961;
            end
    9670  : begin
              real_value= -22395;
              imag_value=23911;
            end
    9671  : begin
              real_value= -26784;
              imag_value=18863;
            end
    9672  : begin
              real_value= -30057;
              imag_value=13030;
            end
    9673  : begin
              real_value= -32077;
              imag_value=6654;
            end
    9674  : begin
              real_value= -32760;
              imag_value=0;
            end
    9675  : begin
              real_value= -32077;
              imag_value=-6654;
            end
    9676  : begin
              real_value= -30057;
              imag_value=-13030;
            end
    9677  : begin
              real_value= -26784;
              imag_value=-18863;
            end
    9678  : begin
              real_value= -22395;
              imag_value=-23911;
            end
    9679  : begin
              real_value= -17072;
              imag_value=-27961;
            end
    9680  : begin
              real_value= -11036;
              imag_value=-30846;
            end
    9681  : begin
              real_value= -4540;
              imag_value=-32445;
            end
    9682  : begin
              real_value= 2142;
              imag_value=-32691;
            end
    9683  : begin
              real_value= 8737;
              imag_value=-31575;
            end
    9684  : begin
              real_value= 14968;
              imag_value=-29142;
            end
    9685  : begin
              real_value= 20575;
              imag_value=-25494;
            end
    9686  : begin
              real_value= 25324;
              imag_value=-20783;
            end
    9687  : begin
              real_value= 29017;
              imag_value=-15206;
            end
    9688  : begin
              real_value= 31501;
              imag_value=-8995;
            end
    9689  : begin
              real_value= 32673;
              imag_value=-2408;
            end
    9690  : begin
              real_value= 32481;
              imag_value=4275;
            end
    9691  : begin
              real_value= 30935;
              imag_value=10783;
            end
    9692  : begin
              real_value= 28100;
              imag_value=16842;
            end
    9693  : begin
              real_value= 24092;
              imag_value=22199;
            end
    9694  : begin
              real_value= 19081;
              imag_value=26630;
            end
    9695  : begin
              real_value= 13274;
              imag_value=29950;
            end
    9696  : begin
              real_value= 6915;
              imag_value=32022;
            end
    9697  : begin
              real_value= 267;
              imag_value=32759;
            end
    9698  : begin
              real_value= -6390;
              imag_value=32131;
            end
    9699  : begin
              real_value= -12784;
              imag_value=30163;
            end
    9700  : begin
              real_value= -18644;
              imag_value=26938;
            end
    9701  : begin
              real_value= -23726;
              imag_value=22589;
            end
    9702  : begin
              real_value= -27820;
              imag_value=17299;
            end
    9703  : begin
              real_value= -30755;
              imag_value=11289;
            end
    9704  : begin
              real_value= -32407;
              imag_value=4806;
            end
    9705  : begin
              real_value= -32707;
              imag_value=-1874;
            end
    9706  : begin
              real_value= -31645;
              imag_value=-8477;
            end
    9707  : begin
              real_value= -29263;
              imag_value=-14728;
            end
    9708  : begin
              real_value= -25661;
              imag_value=-20365;
            end
    9709  : begin
              real_value= -20988;
              imag_value=-25154;
            end
    9710  : begin
              real_value= -15442;
              imag_value=-28892;
            end
    9711  : begin
              real_value= -9253;
              imag_value=-31426;
            end
    9712  : begin
              real_value= -2676;
              imag_value=-32651;
            end
    9713  : begin
              real_value= 4009;
              imag_value=-32515;
            end
    9714  : begin
              real_value= 10529;
              imag_value=-31023;
            end
    9715  : begin
              real_value= 16611;
              imag_value=-28236;
            end
    9716  : begin
              real_value= 22001;
              imag_value=-24274;
            end
    9717  : begin
              real_value= 26472;
              imag_value=-19299;
            end
    9718  : begin
              real_value= 29841;
              imag_value=-13520;
            end
    9719  : begin
              real_value= 31965;
              imag_value=-7177;
            end
    9720  : begin
              real_value= 32757;
              imag_value=-535;
            end
    9721  : begin
              real_value= 32183;
              imag_value=6127;
            end
    9722  : begin
              real_value= 30267;
              imag_value=12537;
            end
    9723  : begin
              real_value= 27090;
              imag_value=18423;
            end
    9724  : begin
              real_value= 22782;
              imag_value=23541;
            end
    9725  : begin
              real_value= 17525;
              imag_value=27678;
            end
    9726  : begin
              real_value= 11539;
              imag_value=30661;
            end
    9727  : begin
              real_value= 5071;
              imag_value=32365;
            end
    9728  : begin
              real_value= -1606;
              imag_value=32721;
            end
    9729  : begin
              real_value= -8219;
              imag_value=31713;
            end
    9730  : begin
              real_value= -14489;
              imag_value=29382;
            end
    9731  : begin
              real_value= -20154;
              imag_value=25826;
            end
    9732  : begin
              real_value= -24981;
              imag_value=21194;
            end
    9733  : begin
              real_value= -28766;
              imag_value=15678;
            end
    9734  : begin
              real_value= -31351;
              imag_value=9508;
            end
    9735  : begin
              real_value= -32629;
              imag_value=2942;
            end
    9736  : begin
              real_value= -32547;
              imag_value=-3742;
            end
    9737  : begin
              real_value= -31107;
              imag_value=-10275;
            end
    9738  : begin
              real_value= -28371;
              imag_value=-16380;
            end
    9739  : begin
              real_value= -24453;
              imag_value=-21801;
            end
    9740  : begin
              real_value= -19515;
              imag_value=-26314;
            end
    9741  : begin
              real_value= -13764;
              imag_value=-29729;
            end
    9742  : begin
              real_value= -7438;
              imag_value=-31905;
            end
    9743  : begin
              real_value= -802;
              imag_value=-32750;
            end
    9744  : begin
              real_value= 5864;
              imag_value=-32231;
            end
    9745  : begin
              real_value= 12288;
              imag_value=-30369;
            end
    9746  : begin
              real_value= 18200;
              imag_value=-27240;
            end
    9747  : begin
              real_value= 23354;
              imag_value=-22974;
            end
    9748  : begin
              real_value= 27534;
              imag_value=-17752;
            end
    9749  : begin
              real_value= 30565;
              imag_value=-11790;
            end
    9750  : begin
              real_value= 32323;
              imag_value=-5336;
            end
    9751  : begin
              real_value= 32733;
              imag_value=1338;
            end
    9752  : begin
              real_value= 31779;
              imag_value=7959;
            end
    9753  : begin
              real_value= 29499;
              imag_value=14248;
            end
    9754  : begin
              real_value= 25990;
              imag_value=19943;
            end
    9755  : begin
              real_value= 21399;
              imag_value=24806;
            end
    9756  : begin
              real_value= 15914;
              imag_value=28636;
            end
    9757  : begin
              real_value= 9765;
              imag_value=31271;
            end
    9758  : begin
              real_value= 3210;
              imag_value=32603;
            end
    9759  : begin
              real_value= -3476;
              imag_value=32575;
            end
    9760  : begin
              real_value= -10021;
              imag_value=31191;
            end
    9761  : begin
              real_value= -16148;
              imag_value=28506;
            end
    9762  : begin
              real_value= -21600;
              imag_value=24630;
            end
    9763  : begin
              real_value= -26152;
              imag_value=19729;
            end
    9764  : begin
              real_value= -29615;
              imag_value=14006;
            end
    9765  : begin
              real_value= -31843;
              imag_value=7699;
            end
    9766  : begin
              real_value= -32743;
              imag_value=1070;
            end
    9767  : begin
              real_value= -32278;
              imag_value=-5599;
            end
    9768  : begin
              real_value= -30468;
              imag_value=-12039;
            end
    9769  : begin
              real_value= -27387;
              imag_value=-17977;
            end
    9770  : begin
              real_value= -23165;
              imag_value=-23165;
            end
    9771  : begin
              real_value= -17977;
              imag_value=-27387;
            end
    9772  : begin
              real_value= -12039;
              imag_value=-30468;
            end
    9773  : begin
              real_value= -5599;
              imag_value=-32278;
            end
    9774  : begin
              real_value= 1070;
              imag_value=-32743;
            end
    9775  : begin
              real_value= 7699;
              imag_value=-31843;
            end
    9776  : begin
              real_value= 14006;
              imag_value=-29615;
            end
    9777  : begin
              real_value= 19729;
              imag_value=-26152;
            end
    9778  : begin
              real_value= 24630;
              imag_value=-21600;
            end
    9779  : begin
              real_value= 28506;
              imag_value=-16148;
            end
    9780  : begin
              real_value= 31191;
              imag_value=-10021;
            end
    9781  : begin
              real_value= 32575;
              imag_value=-3476;
            end
    9782  : begin
              real_value= 32603;
              imag_value=3210;
            end
    9783  : begin
              real_value= 31271;
              imag_value=9765;
            end
    9784  : begin
              real_value= 28636;
              imag_value=15914;
            end
    9785  : begin
              real_value= 24806;
              imag_value=21399;
            end
    9786  : begin
              real_value= 19943;
              imag_value=25990;
            end
    9787  : begin
              real_value= 14248;
              imag_value=29499;
            end
    9788  : begin
              real_value= 7959;
              imag_value=31779;
            end
    9789  : begin
              real_value= 1338;
              imag_value=32733;
            end
    9790  : begin
              real_value= -5336;
              imag_value=32323;
            end
    9791  : begin
              real_value= -11790;
              imag_value=30565;
            end
    9792  : begin
              real_value= -17752;
              imag_value=27534;
            end
    9793  : begin
              real_value= -22974;
              imag_value=23354;
            end
    9794  : begin
              real_value= -27240;
              imag_value=18200;
            end
    9795  : begin
              real_value= -30369;
              imag_value=12288;
            end
    9796  : begin
              real_value= -32231;
              imag_value=5864;
            end
    9797  : begin
              real_value= -32750;
              imag_value=-802;
            end
    9798  : begin
              real_value= -31905;
              imag_value=-7438;
            end
    9799  : begin
              real_value= -29729;
              imag_value=-13764;
            end
    9800  : begin
              real_value= -26314;
              imag_value=-19515;
            end
    9801  : begin
              real_value= -21801;
              imag_value=-24453;
            end
    9802  : begin
              real_value= -16380;
              imag_value=-28371;
            end
    9803  : begin
              real_value= -10275;
              imag_value=-31107;
            end
    9804  : begin
              real_value= -3742;
              imag_value=-32547;
            end
    9805  : begin
              real_value= 2942;
              imag_value=-32629;
            end
    9806  : begin
              real_value= 9508;
              imag_value=-31351;
            end
    9807  : begin
              real_value= 15678;
              imag_value=-28766;
            end
    9808  : begin
              real_value= 21194;
              imag_value=-24981;
            end
    9809  : begin
              real_value= 25826;
              imag_value=-20154;
            end
    9810  : begin
              real_value= 29382;
              imag_value=-14489;
            end
    9811  : begin
              real_value= 31713;
              imag_value=-8219;
            end
    9812  : begin
              real_value= 32721;
              imag_value=-1606;
            end
    9813  : begin
              real_value= 32365;
              imag_value=5071;
            end
    9814  : begin
              real_value= 30661;
              imag_value=11539;
            end
    9815  : begin
              real_value= 27678;
              imag_value=17525;
            end
    9816  : begin
              real_value= 23541;
              imag_value=22782;
            end
    9817  : begin
              real_value= 18423;
              imag_value=27090;
            end
    9818  : begin
              real_value= 12537;
              imag_value=30267;
            end
    9819  : begin
              real_value= 6127;
              imag_value=32183;
            end
    9820  : begin
              real_value= -535;
              imag_value=32757;
            end
    9821  : begin
              real_value= -7177;
              imag_value=31965;
            end
    9822  : begin
              real_value= -13520;
              imag_value=29841;
            end
    9823  : begin
              real_value= -19299;
              imag_value=26472;
            end
    9824  : begin
              real_value= -24274;
              imag_value=22001;
            end
    9825  : begin
              real_value= -28236;
              imag_value=16611;
            end
    9826  : begin
              real_value= -31023;
              imag_value=10529;
            end
    9827  : begin
              real_value= -32515;
              imag_value=4009;
            end
    9828  : begin
              real_value= -32651;
              imag_value=-2676;
            end
    9829  : begin
              real_value= -31426;
              imag_value=-9253;
            end
    9830  : begin
              real_value= -28892;
              imag_value=-15442;
            end
    9831  : begin
              real_value= -25154;
              imag_value=-20988;
            end
    9832  : begin
              real_value= -20365;
              imag_value=-25661;
            end
    9833  : begin
              real_value= -14728;
              imag_value=-29263;
            end
    9834  : begin
              real_value= -8477;
              imag_value=-31645;
            end
    9835  : begin
              real_value= -1874;
              imag_value=-32707;
            end
    9836  : begin
              real_value= 4806;
              imag_value=-32407;
            end
    9837  : begin
              real_value= 11289;
              imag_value=-30755;
            end
    9838  : begin
              real_value= 17299;
              imag_value=-27820;
            end
    9839  : begin
              real_value= 22589;
              imag_value=-23726;
            end
    9840  : begin
              real_value= 26938;
              imag_value=-18644;
            end
    9841  : begin
              real_value= 30163;
              imag_value=-12784;
            end
    9842  : begin
              real_value= 32131;
              imag_value=-6390;
            end
    9843  : begin
              real_value= 32759;
              imag_value=267;
            end
    9844  : begin
              real_value= 32022;
              imag_value=6915;
            end
    9845  : begin
              real_value= 29950;
              imag_value=13274;
            end
    9846  : begin
              real_value= 26630;
              imag_value=19081;
            end
    9847  : begin
              real_value= 22199;
              imag_value=24092;
            end
    9848  : begin
              real_value= 16842;
              imag_value=28100;
            end
    9849  : begin
              real_value= 10783;
              imag_value=30935;
            end
    9850  : begin
              real_value= 4275;
              imag_value=32481;
            end
    9851  : begin
              real_value= -2408;
              imag_value=32673;
            end
    9852  : begin
              real_value= -8995;
              imag_value=31501;
            end
    9853  : begin
              real_value= -15206;
              imag_value=29017;
            end
    9854  : begin
              real_value= -20783;
              imag_value=25324;
            end
    9855  : begin
              real_value= -25494;
              imag_value=20575;
            end
    9856  : begin
              real_value= -29142;
              imag_value=14968;
            end
    9857  : begin
              real_value= -31575;
              imag_value=8737;
            end
    9858  : begin
              real_value= -32691;
              imag_value=2142;
            end
    9859  : begin
              real_value= -32445;
              imag_value=-4540;
            end
    9860  : begin
              real_value= -30846;
              imag_value=-11036;
            end
    9861  : begin
              real_value= -27961;
              imag_value=-17072;
            end
    9862  : begin
              real_value= -23911;
              imag_value=-22395;
            end
    9863  : begin
              real_value= -18863;
              imag_value=-26784;
            end
    9864  : begin
              real_value= -13030;
              imag_value=-30057;
            end
    9865  : begin
              real_value= -6654;
              imag_value=-32077;
            end
    9866  : begin
              real_value= 0;
              imag_value=-32760;
            end
    9867  : begin
              real_value= 6654;
              imag_value=-32077;
            end
    9868  : begin
              real_value= 13030;
              imag_value=-30057;
            end
    9869  : begin
              real_value= 18863;
              imag_value=-26784;
            end
    9870  : begin
              real_value= 23911;
              imag_value=-22395;
            end
    9871  : begin
              real_value= 27961;
              imag_value=-17072;
            end
    9872  : begin
              real_value= 30846;
              imag_value=-11036;
            end
    9873  : begin
              real_value= 32445;
              imag_value=-4540;
            end
    9874  : begin
              real_value= 32691;
              imag_value=2142;
            end
    9875  : begin
              real_value= 31575;
              imag_value=8737;
            end
    9876  : begin
              real_value= 29142;
              imag_value=14968;
            end
    9877  : begin
              real_value= 25494;
              imag_value=20575;
            end
    9878  : begin
              real_value= 20783;
              imag_value=25324;
            end
    9879  : begin
              real_value= 15206;
              imag_value=29017;
            end
    9880  : begin
              real_value= 8995;
              imag_value=31501;
            end
    9881  : begin
              real_value= 2408;
              imag_value=32673;
            end
    9882  : begin
              real_value= -4275;
              imag_value=32481;
            end
    9883  : begin
              real_value= -10783;
              imag_value=30935;
            end
    9884  : begin
              real_value= -16842;
              imag_value=28100;
            end
    9885  : begin
              real_value= -22199;
              imag_value=24092;
            end
    9886  : begin
              real_value= -26630;
              imag_value=19081;
            end
    9887  : begin
              real_value= -29950;
              imag_value=13274;
            end
    9888  : begin
              real_value= -32022;
              imag_value=6915;
            end
    9889  : begin
              real_value= -32759;
              imag_value=267;
            end
    9890  : begin
              real_value= -32131;
              imag_value=-6390;
            end
    9891  : begin
              real_value= -30163;
              imag_value=-12784;
            end
    9892  : begin
              real_value= -26938;
              imag_value=-18644;
            end
    9893  : begin
              real_value= -22589;
              imag_value=-23726;
            end
    9894  : begin
              real_value= -17299;
              imag_value=-27820;
            end
    9895  : begin
              real_value= -11289;
              imag_value=-30755;
            end
    9896  : begin
              real_value= -4806;
              imag_value=-32407;
            end
    9897  : begin
              real_value= 1874;
              imag_value=-32707;
            end
    9898  : begin
              real_value= 8477;
              imag_value=-31645;
            end
    9899  : begin
              real_value= 14728;
              imag_value=-29263;
            end
    9900  : begin
              real_value= 20365;
              imag_value=-25661;
            end
    9901  : begin
              real_value= 25154;
              imag_value=-20988;
            end
    9902  : begin
              real_value= 28892;
              imag_value=-15442;
            end
    9903  : begin
              real_value= 31426;
              imag_value=-9253;
            end
    9904  : begin
              real_value= 32651;
              imag_value=-2676;
            end
    9905  : begin
              real_value= 32515;
              imag_value=4009;
            end
    9906  : begin
              real_value= 31023;
              imag_value=10529;
            end
    9907  : begin
              real_value= 28236;
              imag_value=16611;
            end
    9908  : begin
              real_value= 24274;
              imag_value=22001;
            end
    9909  : begin
              real_value= 19299;
              imag_value=26472;
            end
    9910  : begin
              real_value= 13520;
              imag_value=29841;
            end
    9911  : begin
              real_value= 7177;
              imag_value=31965;
            end
    9912  : begin
              real_value= 535;
              imag_value=32757;
            end
    9913  : begin
              real_value= -6127;
              imag_value=32183;
            end
    9914  : begin
              real_value= -12537;
              imag_value=30267;
            end
    9915  : begin
              real_value= -18423;
              imag_value=27090;
            end
    9916  : begin
              real_value= -23541;
              imag_value=22782;
            end
    9917  : begin
              real_value= -27678;
              imag_value=17525;
            end
    9918  : begin
              real_value= -30661;
              imag_value=11539;
            end
    9919  : begin
              real_value= -32365;
              imag_value=5071;
            end
    9920  : begin
              real_value= -32721;
              imag_value=-1606;
            end
    9921  : begin
              real_value= -31713;
              imag_value=-8219;
            end
    9922  : begin
              real_value= -29382;
              imag_value=-14489;
            end
    9923  : begin
              real_value= -25826;
              imag_value=-20154;
            end
    9924  : begin
              real_value= -21194;
              imag_value=-24981;
            end
    9925  : begin
              real_value= -15678;
              imag_value=-28766;
            end
    9926  : begin
              real_value= -9508;
              imag_value=-31351;
            end
    9927  : begin
              real_value= -2942;
              imag_value=-32629;
            end
    9928  : begin
              real_value= 3742;
              imag_value=-32547;
            end
    9929  : begin
              real_value= 10275;
              imag_value=-31107;
            end
    9930  : begin
              real_value= 16380;
              imag_value=-28371;
            end
    9931  : begin
              real_value= 21801;
              imag_value=-24453;
            end
    9932  : begin
              real_value= 26314;
              imag_value=-19515;
            end
    9933  : begin
              real_value= 29729;
              imag_value=-13764;
            end
    9934  : begin
              real_value= 31905;
              imag_value=-7438;
            end
    9935  : begin
              real_value= 32750;
              imag_value=-802;
            end
    9936  : begin
              real_value= 32231;
              imag_value=5864;
            end
    9937  : begin
              real_value= 30369;
              imag_value=12288;
            end
    9938  : begin
              real_value= 27240;
              imag_value=18200;
            end
    9939  : begin
              real_value= 22974;
              imag_value=23354;
            end
    9940  : begin
              real_value= 17752;
              imag_value=27534;
            end
    9941  : begin
              real_value= 11790;
              imag_value=30565;
            end
    9942  : begin
              real_value= 5336;
              imag_value=32323;
            end
    9943  : begin
              real_value= -1338;
              imag_value=32733;
            end
    9944  : begin
              real_value= -7959;
              imag_value=31779;
            end
    9945  : begin
              real_value= -14248;
              imag_value=29499;
            end
    9946  : begin
              real_value= -19943;
              imag_value=25990;
            end
    9947  : begin
              real_value= -24806;
              imag_value=21399;
            end
    9948  : begin
              real_value= -28636;
              imag_value=15914;
            end
    9949  : begin
              real_value= -31271;
              imag_value=9765;
            end
    9950  : begin
              real_value= -32603;
              imag_value=3210;
            end
    9951  : begin
              real_value= -32575;
              imag_value=-3476;
            end
    9952  : begin
              real_value= -31191;
              imag_value=-10021;
            end
    9953  : begin
              real_value= -28506;
              imag_value=-16148;
            end
    9954  : begin
              real_value= -24630;
              imag_value=-21600;
            end
    9955  : begin
              real_value= -19729;
              imag_value=-26152;
            end
    9956  : begin
              real_value= -14006;
              imag_value=-29615;
            end
    9957  : begin
              real_value= -7699;
              imag_value=-31843;
            end
    9958  : begin
              real_value= -1070;
              imag_value=-32743;
            end
    9959  : begin
              real_value= 5599;
              imag_value=-32278;
            end
    9960  : begin
              real_value= 12039;
              imag_value=-30468;
            end
    9961  : begin
              real_value= 17977;
              imag_value=-27387;
            end
    9962  : begin
              real_value= 23165;
              imag_value=-23165;
            end
    9963  : begin
              real_value= 27387;
              imag_value=-17977;
            end
    9964  : begin
              real_value= 30468;
              imag_value=-12039;
            end
    9965  : begin
              real_value= 32278;
              imag_value=-5599;
            end
    9966  : begin
              real_value= 32743;
              imag_value=1070;
            end
    9967  : begin
              real_value= 31843;
              imag_value=7699;
            end
    9968  : begin
              real_value= 29615;
              imag_value=14006;
            end
    9969  : begin
              real_value= 26152;
              imag_value=19729;
            end
    9970  : begin
              real_value= 21600;
              imag_value=24630;
            end
    9971  : begin
              real_value= 16148;
              imag_value=28506;
            end
    9972  : begin
              real_value= 10021;
              imag_value=31191;
            end
    9973  : begin
              real_value= 3476;
              imag_value=32575;
            end
    9974  : begin
              real_value= -3210;
              imag_value=32603;
            end
    9975  : begin
              real_value= -9765;
              imag_value=31271;
            end
    9976  : begin
              real_value= -15914;
              imag_value=28636;
            end
    9977  : begin
              real_value= -21399;
              imag_value=24806;
            end
    9978  : begin
              real_value= -25990;
              imag_value=19943;
            end
    9979  : begin
              real_value= -29499;
              imag_value=14248;
            end
    9980  : begin
              real_value= -31779;
              imag_value=7959;
            end
    9981  : begin
              real_value= -32733;
              imag_value=1338;
            end
    9982  : begin
              real_value= -32323;
              imag_value=-5336;
            end
    9983  : begin
              real_value= -30565;
              imag_value=-11790;
            end
    9984  : begin
              real_value= -27534;
              imag_value=-17752;
            end
    9985  : begin
              real_value= -23354;
              imag_value=-22974;
            end
    9986  : begin
              real_value= -18200;
              imag_value=-27240;
            end
    9987  : begin
              real_value= -12288;
              imag_value=-30369;
            end
    9988  : begin
              real_value= -5864;
              imag_value=-32231;
            end
    9989  : begin
              real_value= 802;
              imag_value=-32750;
            end
    9990  : begin
              real_value= 7438;
              imag_value=-31905;
            end
    9991  : begin
              real_value= 13764;
              imag_value=-29729;
            end
    9992  : begin
              real_value= 19515;
              imag_value=-26314;
            end
    9993  : begin
              real_value= 24453;
              imag_value=-21801;
            end
    9994  : begin
              real_value= 28371;
              imag_value=-16380;
            end
    9995  : begin
              real_value= 31107;
              imag_value=-10275;
            end
    9996  : begin
              real_value= 32547;
              imag_value=-3742;
            end
    9997  : begin
              real_value= 32629;
              imag_value=2942;
            end
    9998  : begin
              real_value= 31351;
              imag_value=9508;
            end
    9999  : begin
              real_value= 28766;
              imag_value=15678;
            end
    10000  : begin
              real_value= 24981;
              imag_value=21194;
            end
    10001 : begin
              real_value= 20154;
              imag_value=25826;
            end
    10002 : begin
              real_value= 14489;
              imag_value=29382;
            end
    10003 : begin
              real_value= 8219;
              imag_value=31713;
            end
    10004 : begin
              real_value= 1606;
              imag_value=32721;
            end
    10005 : begin
              real_value= -5071;
              imag_value=32365;
            end
    10006 : begin
              real_value= -11539;
              imag_value=30661;
            end
    10007 : begin
              real_value= -17525;
              imag_value=27678;
            end
    10008 : begin
              real_value= -22782;
              imag_value=23541;
            end
    10009 : begin
              real_value= -27090;
              imag_value=18423;
            end
    10010 : begin
              real_value= -30267;
              imag_value=12537;
            end
    10011 : begin
              real_value= -32183;
              imag_value=6127;
            end
    10012 : begin
              real_value= -32757;
              imag_value=-535;
            end
    10013 : begin
              real_value= -31965;
              imag_value=-7177;
            end
    10014 : begin
              real_value= -29841;
              imag_value=-13520;
            end
    10015 : begin
              real_value= -26472;
              imag_value=-19299;
            end
    10016 : begin
              real_value= -22001;
              imag_value=-24274;
            end
    10017 : begin
              real_value= -16611;
              imag_value=-28236;
            end
    10018 : begin
              real_value= -10529;
              imag_value=-31023;
            end
    10019 : begin
              real_value= -4009;
              imag_value=-32515;
            end
    10020 : begin
              real_value= 2676;
              imag_value=-32651;
            end
    10021 : begin
              real_value= 9253;
              imag_value=-31426;
            end
    10022 : begin
              real_value= 15442;
              imag_value=-28892;
            end
    10023 : begin
              real_value= 20988;
              imag_value=-25154;
            end
    10024 : begin
              real_value= 25661;
              imag_value=-20365;
            end
    10025 : begin
              real_value= 29263;
              imag_value=-14728;
            end
    10026 : begin
              real_value= 31645;
              imag_value=-8477;
            end
    10027 : begin
              real_value= 32707;
              imag_value=-1874;
            end
    10028 : begin
              real_value= 32407;
              imag_value=4806;
            end
    10029 : begin
              real_value= 30755;
              imag_value=11289;
            end
    10030 : begin
              real_value= 27820;
              imag_value=17299;
            end
    10031 : begin
              real_value= 23726;
              imag_value=22589;
            end
    10032 : begin
              real_value= 18644;
              imag_value=26938;
            end
    10033 : begin
              real_value= 12784;
              imag_value=30163;
            end
    10034 : begin
              real_value= 6390;
              imag_value=32131;
            end
    10035 : begin
              real_value= -267;
              imag_value=32759;
            end
    10036 : begin
              real_value= -6915;
              imag_value=32022;
            end
    10037 : begin
              real_value= -13274;
              imag_value=29950;
            end
    10038 : begin
              real_value= -19081;
              imag_value=26630;
            end
    10039 : begin
              real_value= -24092;
              imag_value=22199;
            end
    10040 : begin
              real_value= -28100;
              imag_value=16842;
            end
    10041 : begin
              real_value= -30935;
              imag_value=10783;
            end
    10042 : begin
              real_value= -32481;
              imag_value=4275;
            end
    10043 : begin
              real_value= -32673;
              imag_value=-2408;
            end
    10044 : begin
              real_value= -31501;
              imag_value=-8995;
            end
    10045 : begin
              real_value= -29017;
              imag_value=-15206;
            end
    10046 : begin
              real_value= -25324;
              imag_value=-20783;
            end
    10047 : begin
              real_value= -20575;
              imag_value=-25494;
            end
    10048 : begin
              real_value= -14968;
              imag_value=-29142;
            end
    10049 : begin
              real_value= -8737;
              imag_value=-31575;
            end
    10050 : begin
              real_value= -2142;
              imag_value=-32691;
            end
    10051 : begin
              real_value= 4540;
              imag_value=-32445;
            end
    10052 : begin
              real_value= 11036;
              imag_value=-30846;
            end
    10053 : begin
              real_value= 17072;
              imag_value=-27961;
            end
    10054 : begin
              real_value= 22395;
              imag_value=-23911;
            end
    10055 : begin
              real_value= 26784;
              imag_value=-18863;
            end
    10056 : begin
              real_value= 30057;
              imag_value=-13030;
            end
    10057 : begin
              real_value= 32077;
              imag_value=-6654;
            end
    10058 : begin
              real_value= 32760;
              imag_value=0;
            end
    10059 : begin
              real_value= 32077;
              imag_value=6654;
            end
    10060 : begin
              real_value= 30057;
              imag_value=13030;
            end
    10061 : begin
              real_value= 26784;
              imag_value=18863;
            end
    10062 : begin
              real_value= 22395;
              imag_value=23911;
            end
    10063 : begin
              real_value= 17072;
              imag_value=27961;
            end
    10064 : begin
              real_value= 11036;
              imag_value=30846;
            end
    10065 : begin
              real_value= 4540;
              imag_value=32445;
            end
    10066 : begin
              real_value= -2142;
              imag_value=32691;
            end
    10067 : begin
              real_value= -8737;
              imag_value=31575;
            end
    10068 : begin
              real_value= -14968;
              imag_value=29142;
            end
    10069 : begin
              real_value= -20575;
              imag_value=25494;
            end
    10070 : begin
              real_value= -25324;
              imag_value=20783;
            end
    10071 : begin
              real_value= -29017;
              imag_value=15206;
            end
    10072 : begin
              real_value= -31501;
              imag_value=8995;
            end
    10073 : begin
              real_value= -32673;
              imag_value=2408;
            end
    10074 : begin
              real_value= -32481;
              imag_value=-4275;
            end
    10075 : begin
              real_value= -30935;
              imag_value=-10783;
            end
    10076 : begin
              real_value= -28100;
              imag_value=-16842;
            end
    10077 : begin
              real_value= -24092;
              imag_value=-22199;
            end
    10078 : begin
              real_value= -19081;
              imag_value=-26630;
            end
    10079 : begin
              real_value= -13274;
              imag_value=-29950;
            end
    10080 : begin
              real_value= -6915;
              imag_value=-32022;
            end
    10081 : begin
              real_value= -267;
              imag_value=-32759;
            end
    10082 : begin
              real_value= 6390;
              imag_value=-32131;
            end
    10083 : begin
              real_value= 12784;
              imag_value=-30163;
            end
    10084 : begin
              real_value= 18644;
              imag_value=-26938;
            end
    10085 : begin
              real_value= 23726;
              imag_value=-22589;
            end
    10086 : begin
              real_value= 27820;
              imag_value=-17299;
            end
    10087 : begin
              real_value= 30755;
              imag_value=-11289;
            end
    10088 : begin
              real_value= 32407;
              imag_value=-4806;
            end
    10089 : begin
              real_value= 32707;
              imag_value=1874;
            end
    10090 : begin
              real_value= 31645;
              imag_value=8477;
            end
    10091 : begin
              real_value= 29263;
              imag_value=14728;
            end
    10092 : begin
              real_value= 25661;
              imag_value=20365;
            end
    10093 : begin
              real_value= 20988;
              imag_value=25154;
            end
    10094 : begin
              real_value= 15442;
              imag_value=28892;
            end
    10095 : begin
              real_value= 9253;
              imag_value=31426;
            end
    10096 : begin
              real_value= 2676;
              imag_value=32651;
            end
    10097 : begin
              real_value= -4009;
              imag_value=32515;
            end
    10098 : begin
              real_value= -10529;
              imag_value=31023;
            end
    10099 : begin
              real_value= -16611;
              imag_value=28236;
            end
    10100 : begin
              real_value= -22001;
              imag_value=24274;
            end
    10101 : begin
              real_value= -26472;
              imag_value=19299;
            end
    10102 : begin
              real_value= -29841;
              imag_value=13520;
            end
    10103 : begin
              real_value= -31965;
              imag_value=7177;
            end
    10104 : begin
              real_value= -32757;
              imag_value=535;
            end
    10105 : begin
              real_value= -32183;
              imag_value=-6127;
            end
    10106 : begin
              real_value= -30267;
              imag_value=-12537;
            end
    10107 : begin
              real_value= -27090;
              imag_value=-18423;
            end
    10108 : begin
              real_value= -22782;
              imag_value=-23541;
            end
    10109 : begin
              real_value= -17525;
              imag_value=-27678;
            end
    10110 : begin
              real_value= -11539;
              imag_value=-30661;
            end
    10111 : begin
              real_value= -5071;
              imag_value=-32365;
            end
    10112 : begin
              real_value= 1606;
              imag_value=-32721;
            end
    10113 : begin
              real_value= 8219;
              imag_value=-31713;
            end
    10114 : begin
              real_value= 14489;
              imag_value=-29382;
            end
    10115 : begin
              real_value= 20154;
              imag_value=-25826;
            end
    10116 : begin
              real_value= 24981;
              imag_value=-21194;
            end
    10117 : begin
              real_value= 28766;
              imag_value=-15678;
            end
    10118 : begin
              real_value= 31351;
              imag_value=-9508;
            end
    10119 : begin
              real_value= 32629;
              imag_value=-2942;
            end
    10120 : begin
              real_value= 32547;
              imag_value=3742;
            end
    10121 : begin
              real_value= 31107;
              imag_value=10275;
            end
    10122 : begin
              real_value= 28371;
              imag_value=16380;
            end
    10123 : begin
              real_value= 24453;
              imag_value=21801;
            end
    10124 : begin
              real_value= 19515;
              imag_value=26314;
            end
    10125 : begin
              real_value= 13764;
              imag_value=29729;
            end
    10126 : begin
              real_value= 7438;
              imag_value=31905;
            end
    10127 : begin
              real_value= 802;
              imag_value=32750;
            end
    10128 : begin
              real_value= -5864;
              imag_value=32231;
            end
    10129 : begin
              real_value= -12288;
              imag_value=30369;
            end
    10130 : begin
              real_value= -18200;
              imag_value=27240;
            end
    10131 : begin
              real_value= -23354;
              imag_value=22974;
            end
    10132 : begin
              real_value= -27534;
              imag_value=17752;
            end
    10133 : begin
              real_value= -30565;
              imag_value=11790;
            end
    10134 : begin
              real_value= -32323;
              imag_value=5336;
            end
    10135 : begin
              real_value= -32733;
              imag_value=-1338;
            end
    10136 : begin
              real_value= -31779;
              imag_value=-7959;
            end
    10137 : begin
              real_value= -29499;
              imag_value=-14248;
            end
    10138 : begin
              real_value= -25990;
              imag_value=-19943;
            end
    10139 : begin
              real_value= -21399;
              imag_value=-24806;
            end
    10140 : begin
              real_value= -15914;
              imag_value=-28636;
            end
    10141 : begin
              real_value= -9765;
              imag_value=-31271;
            end
    10142 : begin
              real_value= -3210;
              imag_value=-32603;
            end
    10143 : begin
              real_value= 3476;
              imag_value=-32575;
            end
    10144 : begin
              real_value= 10021;
              imag_value=-31191;
            end
    10145 : begin
              real_value= 16148;
              imag_value=-28506;
            end
    10146 : begin
              real_value= 21600;
              imag_value=-24630;
            end
    10147 : begin
              real_value= 26152;
              imag_value=-19729;
            end
    10148 : begin
              real_value= 29615;
              imag_value=-14006;
            end
    10149 : begin
              real_value= 31843;
              imag_value=-7699;
            end
    10150 : begin
              real_value= 32743;
              imag_value=-1070;
            end
    10151 : begin
              real_value= 32278;
              imag_value=5599;
            end
    10152 : begin
              real_value= 30468;
              imag_value=12039;
            end
    10153 : begin
              real_value= 27387;
              imag_value=17977;
            end
    10154 : begin
              real_value= 23165;
              imag_value=23165;
            end
    10155 : begin
              real_value= 17977;
              imag_value=27387;
            end
    10156 : begin
              real_value= 12039;
              imag_value=30468;
            end
    10157 : begin
              real_value= 5599;
              imag_value=32278;
            end
    10158 : begin
              real_value= -1070;
              imag_value=32743;
            end
    10159 : begin
              real_value= -7699;
              imag_value=31843;
            end
    10160 : begin
              real_value= -14006;
              imag_value=29615;
            end
    10161 : begin
              real_value= -19729;
              imag_value=26152;
            end
    10162 : begin
              real_value= -24630;
              imag_value=21600;
            end
    10163 : begin
              real_value= -28506;
              imag_value=16148;
            end
    10164 : begin
              real_value= -31191;
              imag_value=10021;
            end
    10165 : begin
              real_value= -32575;
              imag_value=3476;
            end
    10166 : begin
              real_value= -32603;
              imag_value=-3210;
            end
    10167 : begin
              real_value= -31271;
              imag_value=-9765;
            end
    10168 : begin
              real_value= -28636;
              imag_value=-15914;
            end
    10169 : begin
              real_value= -24806;
              imag_value=-21399;
            end
    10170 : begin
              real_value= -19943;
              imag_value=-25990;
            end
    10171 : begin
              real_value= -14248;
              imag_value=-29499;
            end
    10172 : begin
              real_value= -7959;
              imag_value=-31779;
            end
    10173 : begin
              real_value= -1338;
              imag_value=-32733;
            end
    10174 : begin
              real_value= 5336;
              imag_value=-32323;
            end
    10175 : begin
              real_value= 11790;
              imag_value=-30565;
            end
    10176 : begin
              real_value= 17752;
              imag_value=-27534;
            end
    10177 : begin
              real_value= 22974;
              imag_value=-23354;
            end
    10178 : begin
              real_value= 27240;
              imag_value=-18200;
            end
    10179 : begin
              real_value= 30369;
              imag_value=-12288;
            end
    10180 : begin
              real_value= 32231;
              imag_value=-5864;
            end
    10181 : begin
              real_value= 32750;
              imag_value=802;
            end
    10182 : begin
              real_value= 31905;
              imag_value=7438;
            end
    10183 : begin
              real_value= 29729;
              imag_value=13764;
            end
    10184 : begin
              real_value= 26314;
              imag_value=19515;
            end
    10185 : begin
              real_value= 21801;
              imag_value=24453;
            end
    10186 : begin
              real_value= 16380;
              imag_value=28371;
            end
    10187 : begin
              real_value= 10275;
              imag_value=31107;
            end
    10188 : begin
              real_value= 3742;
              imag_value=32547;
            end
    10189 : begin
              real_value= -2942;
              imag_value=32629;
            end
    10190 : begin
              real_value= -9508;
              imag_value=31351;
            end
    10191 : begin
              real_value= -15678;
              imag_value=28766;
            end
    10192 : begin
              real_value= -21194;
              imag_value=24981;
            end
    10193 : begin
              real_value= -25826;
              imag_value=20154;
            end
    10194 : begin
              real_value= -29382;
              imag_value=14489;
            end
    10195 : begin
              real_value= -31713;
              imag_value=8219;
            end
    10196 : begin
              real_value= -32721;
              imag_value=1606;
            end
    10197 : begin
              real_value= -32365;
              imag_value=-5071;
            end
    10198 : begin
              real_value= -30661;
              imag_value=-11539;
            end
    10199 : begin
              real_value= -27678;
              imag_value=-17525;
            end
    10200 : begin
              real_value= -23541;
              imag_value=-22782;
            end
    10201 : begin
              real_value= -18423;
              imag_value=-27090;
            end
    10202 : begin
              real_value= -12537;
              imag_value=-30267;
            end
    10203 : begin
              real_value= -6127;
              imag_value=-32183;
            end
    10204 : begin
              real_value= 535;
              imag_value=-32757;
            end
    10205 : begin
              real_value= 7177;
              imag_value=-31965;
            end
    10206 : begin
              real_value= 13520;
              imag_value=-29841;
            end
    10207 : begin
              real_value= 19299;
              imag_value=-26472;
            end
    10208 : begin
              real_value= 24274;
              imag_value=-22001;
            end
    10209 : begin
              real_value= 28236;
              imag_value=-16611;
            end
    10210 : begin
              real_value= 31023;
              imag_value=-10529;
            end
    10211 : begin
              real_value= 32515;
              imag_value=-4009;
            end
    10212 : begin
              real_value= 32651;
              imag_value=2676;
            end
    10213 : begin
              real_value= 31426;
              imag_value=9253;
            end
    10214 : begin
              real_value= 28892;
              imag_value=15442;
            end
    10215 : begin
              real_value= 25154;
              imag_value=20988;
            end
    10216 : begin
              real_value= 20365;
              imag_value=25661;
            end
    10217 : begin
              real_value= 14728;
              imag_value=29263;
            end
    10218 : begin
              real_value= 8477;
              imag_value=31645;
            end
    10219 : begin
              real_value= 1874;
              imag_value=32707;
            end
    10220 : begin
              real_value= -4806;
              imag_value=32407;
            end
    10221 : begin
              real_value= -11289;
              imag_value=30755;
            end
    10222 : begin
              real_value= -17299;
              imag_value=27820;
            end
    10223 : begin
              real_value= -22589;
              imag_value=23726;
            end
    10224 : begin
              real_value= -26938;
              imag_value=18644;
            end
    10225 : begin
              real_value= -30163;
              imag_value=12784;
            end
    10226 : begin
              real_value= -32131;
              imag_value=6390;
            end
    10227 : begin
              real_value= -32759;
              imag_value=-267;
            end
    10228 : begin
              real_value= -32022;
              imag_value=-6915;
            end
    10229 : begin
              real_value= -29950;
              imag_value=-13274;
            end
    10230 : begin
              real_value= -26630;
              imag_value=-19081;
            end
    10231 : begin
              real_value= -22199;
              imag_value=-24092;
            end
    10232 : begin
              real_value= -16842;
              imag_value=-28100;
            end
    10233 : begin
              real_value= -10783;
              imag_value=-30935;
            end
    10234 : begin
              real_value= -4275;
              imag_value=-32481;
            end
    10235 : begin
              real_value= 2408;
              imag_value=-32673;
            end
    10236 : begin
              real_value= 8995;
              imag_value=-31501;
            end
    10237 : begin
              real_value= 15206;
              imag_value=-29017;
            end
    10238 : begin
              real_value= 20783;
              imag_value=-25324;
            end
    10239 : begin
              real_value= 25494;
              imag_value=-20575;
            end
    10240 : begin
              real_value= 29142;
              imag_value=-14968;
            end
    10241 : begin
              real_value= 31575;
              imag_value=-8737;
            end
    10242 : begin
              real_value= 32691;
              imag_value=-2142;
            end
    10243 : begin
              real_value= 32445;
              imag_value=4540;
            end
    10244 : begin
              real_value= 30846;
              imag_value=11036;
            end
    10245 : begin
              real_value= 27961;
              imag_value=17072;
            end
    10246 : begin
              real_value= 23911;
              imag_value=22395;
            end
    10247 : begin
              real_value= 18863;
              imag_value=26784;
            end
    10248 : begin
              real_value= 13030;
              imag_value=30057;
            end
    10249 : begin
              real_value= 6654;
              imag_value=32077;
            end
    10250 : begin
              real_value= 0;
              imag_value=32760;
            end
    10251 : begin
              real_value= -6654;
              imag_value=32077;
            end
    10252 : begin
              real_value= -13030;
              imag_value=30057;
            end
    10253 : begin
              real_value= -18863;
              imag_value=26784;
            end
    10254 : begin
              real_value= -23911;
              imag_value=22395;
            end
    10255 : begin
              real_value= -27961;
              imag_value=17072;
            end
    10256 : begin
              real_value= -30846;
              imag_value=11036;
            end
    10257 : begin
              real_value= -32445;
              imag_value=4540;
            end
    10258 : begin
              real_value= -32691;
              imag_value=-2142;
            end
    10259 : begin
              real_value= -31575;
              imag_value=-8737;
            end
    10260 : begin
              real_value= -29142;
              imag_value=-14968;
            end
    10261 : begin
              real_value= -25494;
              imag_value=-20575;
            end
    10262 : begin
              real_value= -20783;
              imag_value=-25324;
            end
    10263 : begin
              real_value= -15206;
              imag_value=-29017;
            end
    10264 : begin
              real_value= -8995;
              imag_value=-31501;
            end
    10265 : begin
              real_value= -2408;
              imag_value=-32673;
            end
    10266 : begin
              real_value= 4275;
              imag_value=-32481;
            end
    10267 : begin
              real_value= 10783;
              imag_value=-30935;
            end
    10268 : begin
              real_value= 16842;
              imag_value=-28100;
            end
    10269 : begin
              real_value= 22199;
              imag_value=-24092;
            end
    10270 : begin
              real_value= 26630;
              imag_value=-19081;
            end
    10271 : begin
              real_value= 29950;
              imag_value=-13274;
            end
    10272 : begin
              real_value= 32022;
              imag_value=-6915;
            end
    10273 : begin
              real_value= 32759;
              imag_value=-267;
            end
    10274 : begin
              real_value= 32131;
              imag_value=6390;
            end
    10275 : begin
              real_value= 30163;
              imag_value=12784;
            end
    10276 : begin
              real_value= 26938;
              imag_value=18644;
            end
    10277 : begin
              real_value= 22589;
              imag_value=23726;
            end
    10278 : begin
              real_value= 17299;
              imag_value=27820;
            end
    10279 : begin
              real_value= 11289;
              imag_value=30755;
            end
    10280 : begin
              real_value= 4806;
              imag_value=32407;
            end
    10281 : begin
              real_value= -1874;
              imag_value=32707;
            end
    10282 : begin
              real_value= -8477;
              imag_value=31645;
            end
    10283 : begin
              real_value= -14728;
              imag_value=29263;
            end
    10284 : begin
              real_value= -20365;
              imag_value=25661;
            end
    10285 : begin
              real_value= -25154;
              imag_value=20988;
            end
    10286 : begin
              real_value= -28892;
              imag_value=15442;
            end
    10287 : begin
              real_value= -31426;
              imag_value=9253;
            end
    10288 : begin
              real_value= -32651;
              imag_value=2676;
            end
    10289 : begin
              real_value= -32515;
              imag_value=-4009;
            end
    10290 : begin
              real_value= -31023;
              imag_value=-10529;
            end
    10291 : begin
              real_value= -28236;
              imag_value=-16611;
            end
    10292 : begin
              real_value= -24274;
              imag_value=-22001;
            end
    10293 : begin
              real_value= -19299;
              imag_value=-26472;
            end
    10294 : begin
              real_value= -13520;
              imag_value=-29841;
            end
    10295 : begin
              real_value= -7177;
              imag_value=-31965;
            end
    10296 : begin
              real_value= -535;
              imag_value=-32757;
            end
    10297 : begin
              real_value= 6127;
              imag_value=-32183;
            end
    10298 : begin
              real_value= 12537;
              imag_value=-30267;
            end
    10299 : begin
              real_value= 18423;
              imag_value=-27090;
            end
    10300 : begin
              real_value= 23541;
              imag_value=-22782;
            end
    10301 : begin
              real_value= 27678;
              imag_value=-17525;
            end
    10302 : begin
              real_value= 30661;
              imag_value=-11539;
            end
    10303 : begin
              real_value= 32365;
              imag_value=-5071;
            end
    10304 : begin
              real_value= 32721;
              imag_value=1606;
            end
    10305 : begin
              real_value= 31713;
              imag_value=8219;
            end
    10306 : begin
              real_value= 29382;
              imag_value=14489;
            end
    10307 : begin
              real_value= 25826;
              imag_value=20154;
            end
    10308 : begin
              real_value= 21194;
              imag_value=24981;
            end
    10309 : begin
              real_value= 15678;
              imag_value=28766;
            end
    10310 : begin
              real_value= 9508;
              imag_value=31351;
            end
    10311 : begin
              real_value= 2942;
              imag_value=32629;
            end
    10312 : begin
              real_value= -3742;
              imag_value=32547;
            end
    10313 : begin
              real_value= -10275;
              imag_value=31107;
            end
    10314 : begin
              real_value= -16380;
              imag_value=28371;
            end
    10315 : begin
              real_value= -21801;
              imag_value=24453;
            end
    10316 : begin
              real_value= -26314;
              imag_value=19515;
            end
    10317 : begin
              real_value= -29729;
              imag_value=13764;
            end
    10318 : begin
              real_value= -31905;
              imag_value=7438;
            end
    10319 : begin
              real_value= -32750;
              imag_value=802;
            end
    10320 : begin
              real_value= -32231;
              imag_value=-5864;
            end
    10321 : begin
              real_value= -30369;
              imag_value=-12288;
            end
    10322 : begin
              real_value= -27240;
              imag_value=-18200;
            end
    10323 : begin
              real_value= -22974;
              imag_value=-23354;
            end
    10324 : begin
              real_value= -17752;
              imag_value=-27534;
            end
    10325 : begin
              real_value= -11790;
              imag_value=-30565;
            end
    10326 : begin
              real_value= -5336;
              imag_value=-32323;
            end
    10327 : begin
              real_value= 1338;
              imag_value=-32733;
            end
    10328 : begin
              real_value= 7959;
              imag_value=-31779;
            end
    10329 : begin
              real_value= 14248;
              imag_value=-29499;
            end
    10330 : begin
              real_value= 19943;
              imag_value=-25990;
            end
    10331 : begin
              real_value= 24806;
              imag_value=-21399;
            end
    10332 : begin
              real_value= 28636;
              imag_value=-15914;
            end
    10333 : begin
              real_value= 31271;
              imag_value=-9765;
            end
    10334 : begin
              real_value= 32603;
              imag_value=-3210;
            end
    10335 : begin
              real_value= 32575;
              imag_value=3476;
            end
    10336 : begin
              real_value= 31191;
              imag_value=10021;
            end
    10337 : begin
              real_value= 28506;
              imag_value=16148;
            end
    10338 : begin
              real_value= 24630;
              imag_value=21600;
            end
    10339 : begin
              real_value= 19729;
              imag_value=26152;
            end
    10340 : begin
              real_value= 14006;
              imag_value=29615;
            end
    10341 : begin
              real_value= 7699;
              imag_value=31843;
            end
    10342 : begin
              real_value= 1070;
              imag_value=32743;
            end
    10343 : begin
              real_value= -5599;
              imag_value=32278;
            end
    10344 : begin
              real_value= -12039;
              imag_value=30468;
            end
    10345 : begin
              real_value= -17977;
              imag_value=27387;
            end
    10346 : begin
              real_value= -23165;
              imag_value=23165;
            end
    10347 : begin
              real_value= -27387;
              imag_value=17977;
            end
    10348 : begin
              real_value= -30468;
              imag_value=12039;
            end
    10349 : begin
              real_value= -32278;
              imag_value=5599;
            end
    10350 : begin
              real_value= -32743;
              imag_value=-1070;
            end
    10351 : begin
              real_value= -31843;
              imag_value=-7699;
            end
    10352 : begin
              real_value= -29615;
              imag_value=-14006;
            end
    10353 : begin
              real_value= -26152;
              imag_value=-19729;
            end
    10354 : begin
              real_value= -21600;
              imag_value=-24630;
            end
    10355 : begin
              real_value= -16148;
              imag_value=-28506;
            end
    10356 : begin
              real_value= -10021;
              imag_value=-31191;
            end
    10357 : begin
              real_value= -3476;
              imag_value=-32575;
            end
    10358 : begin
              real_value= 3210;
              imag_value=-32603;
            end
    10359 : begin
              real_value= 9765;
              imag_value=-31271;
            end
    10360 : begin
              real_value= 15914;
              imag_value=-28636;
            end
    10361 : begin
              real_value= 21399;
              imag_value=-24806;
            end
    10362 : begin
              real_value= 25990;
              imag_value=-19943;
            end
    10363 : begin
              real_value= 29499;
              imag_value=-14248;
            end
    10364 : begin
              real_value= 31779;
              imag_value=-7959;
            end
    10365 : begin
              real_value= 32733;
              imag_value=-1338;
            end
    10366 : begin
              real_value= 32323;
              imag_value=5336;
            end
    10367 : begin
              real_value= 30565;
              imag_value=11790;
            end
    10368 : begin
              real_value= 27534;
              imag_value=17752;
            end
    10369 : begin
              real_value= 23354;
              imag_value=22974;
            end
    10370 : begin
              real_value= 18200;
              imag_value=27240;
            end
    10371 : begin
              real_value= 12288;
              imag_value=30369;
            end
    10372 : begin
              real_value= 5864;
              imag_value=32231;
            end
    10373 : begin
              real_value= -802;
              imag_value=32750;
            end
    10374 : begin
              real_value= -7438;
              imag_value=31905;
            end
    10375 : begin
              real_value= -13764;
              imag_value=29729;
            end
    10376 : begin
              real_value= -19515;
              imag_value=26314;
            end
    10377 : begin
              real_value= -24453;
              imag_value=21801;
            end
    10378 : begin
              real_value= -28371;
              imag_value=16380;
            end
    10379 : begin
              real_value= -31107;
              imag_value=10275;
            end
    10380 : begin
              real_value= -32547;
              imag_value=3742;
            end
    10381 : begin
              real_value= -32629;
              imag_value=-2942;
            end
    10382 : begin
              real_value= -31351;
              imag_value=-9508;
            end
    10383 : begin
              real_value= -28766;
              imag_value=-15678;
            end
    10384 : begin
              real_value= -24981;
              imag_value=-21194;
            end
    10385 : begin
              real_value= -20154;
              imag_value=-25826;
            end
    10386 : begin
              real_value= -14489;
              imag_value=-29382;
            end
    10387 : begin
              real_value= -8219;
              imag_value=-31713;
            end
    10388 : begin
              real_value= -1606;
              imag_value=-32721;
            end
    10389 : begin
              real_value= 5071;
              imag_value=-32365;
            end
    10390 : begin
              real_value= 11539;
              imag_value=-30661;
            end
    10391 : begin
              real_value= 17525;
              imag_value=-27678;
            end
    10392 : begin
              real_value= 22782;
              imag_value=-23541;
            end
    10393 : begin
              real_value= 27090;
              imag_value=-18423;
            end
    10394 : begin
              real_value= 30267;
              imag_value=-12537;
            end
    10395 : begin
              real_value= 32183;
              imag_value=-6127;
            end
    10396 : begin
              real_value= 32757;
              imag_value=535;
            end
    10397 : begin
              real_value= 31965;
              imag_value=7177;
            end
    10398 : begin
              real_value= 29841;
              imag_value=13520;
            end
    10399 : begin
              real_value= 26472;
              imag_value=19299;
            end
    10400 : begin
              real_value= 22001;
              imag_value=24274;
            end
    10401 : begin
              real_value= 16611;
              imag_value=28236;
            end
    10402 : begin
              real_value= 10529;
              imag_value=31023;
            end
    10403 : begin
              real_value= 4009;
              imag_value=32515;
            end
    10404 : begin
              real_value= -2676;
              imag_value=32651;
            end
    10405 : begin
              real_value= -9253;
              imag_value=31426;
            end
    10406 : begin
              real_value= -15442;
              imag_value=28892;
            end
    10407 : begin
              real_value= -20988;
              imag_value=25154;
            end
    10408 : begin
              real_value= -25661;
              imag_value=20365;
            end
    10409 : begin
              real_value= -29263;
              imag_value=14728;
            end
    10410 : begin
              real_value= -31645;
              imag_value=8477;
            end
    10411 : begin
              real_value= -32707;
              imag_value=1874;
            end
    10412 : begin
              real_value= -32407;
              imag_value=-4806;
            end
    10413 : begin
              real_value= -30755;
              imag_value=-11289;
            end
    10414 : begin
              real_value= -27820;
              imag_value=-17299;
            end
    10415 : begin
              real_value= -23726;
              imag_value=-22589;
            end
    10416 : begin
              real_value= -18644;
              imag_value=-26938;
            end
    10417 : begin
              real_value= -12784;
              imag_value=-30163;
            end
    10418 : begin
              real_value= -6390;
              imag_value=-32131;
            end
    10419 : begin
              real_value= 267;
              imag_value=-32759;
            end
    10420 : begin
              real_value= 6915;
              imag_value=-32022;
            end
    10421 : begin
              real_value= 13274;
              imag_value=-29950;
            end
    10422 : begin
              real_value= 19081;
              imag_value=-26630;
            end
    10423 : begin
              real_value= 24092;
              imag_value=-22199;
            end
    10424 : begin
              real_value= 28100;
              imag_value=-16842;
            end
    10425 : begin
              real_value= 30935;
              imag_value=-10783;
            end
    10426 : begin
              real_value= 32481;
              imag_value=-4275;
            end
    10427 : begin
              real_value= 32673;
              imag_value=2408;
            end
    10428 : begin
              real_value= 31501;
              imag_value=8995;
            end
    10429 : begin
              real_value= 29017;
              imag_value=15206;
            end
    10430 : begin
              real_value= 25324;
              imag_value=20783;
            end
    10431 : begin
              real_value= 20575;
              imag_value=25494;
            end
    10432 : begin
              real_value= 14968;
              imag_value=29142;
            end
    10433 : begin
              real_value= 8737;
              imag_value=31575;
            end
    10434 : begin
              real_value= 2142;
              imag_value=32691;
            end
    10435 : begin
              real_value= -4540;
              imag_value=32445;
            end
    10436 : begin
              real_value= -11036;
              imag_value=30846;
            end
    10437 : begin
              real_value= -17072;
              imag_value=27961;
            end
    10438 : begin
              real_value= -22395;
              imag_value=23911;
            end
    10439 : begin
              real_value= -26784;
              imag_value=18863;
            end
    10440 : begin
              real_value= -30057;
              imag_value=13030;
            end
    10441 : begin
              real_value= -32077;
              imag_value=6654;
            end
    10442 : begin
              real_value= -32760;
              imag_value=0;
            end
    10443 : begin
              real_value= -32077;
              imag_value=-6654;
            end
    10444 : begin
              real_value= -30057;
              imag_value=-13030;
            end
    10445 : begin
              real_value= -26784;
              imag_value=-18863;
            end
    10446 : begin
              real_value= -22395;
              imag_value=-23911;
            end
    10447 : begin
              real_value= -17072;
              imag_value=-27961;
            end
    10448 : begin
              real_value= -11036;
              imag_value=-30846;
            end
    10449 : begin
              real_value= -4540;
              imag_value=-32445;
            end
    10450 : begin
              real_value= 2142;
              imag_value=-32691;
            end
    10451 : begin
              real_value= 8737;
              imag_value=-31575;
            end
    10452 : begin
              real_value= 14968;
              imag_value=-29142;
            end
    10453 : begin
              real_value= 20575;
              imag_value=-25494;
            end
    10454 : begin
              real_value= 25324;
              imag_value=-20783;
            end
    10455 : begin
              real_value= 29017;
              imag_value=-15206;
            end
    10456 : begin
              real_value= 31501;
              imag_value=-8995;
            end
    10457 : begin
              real_value= 32673;
              imag_value=-2408;
            end
    10458 : begin
              real_value= 32481;
              imag_value=4275;
            end
    10459 : begin
              real_value= 30935;
              imag_value=10783;
            end
    10460 : begin
              real_value= 28100;
              imag_value=16842;
            end
    10461 : begin
              real_value= 24092;
              imag_value=22199;
            end
    10462 : begin
              real_value= 19081;
              imag_value=26630;
            end
    10463 : begin
              real_value= 13274;
              imag_value=29950;
            end
    10464 : begin
              real_value= 6915;
              imag_value=32022;
            end
    10465 : begin
              real_value= 267;
              imag_value=32759;
            end
    10466 : begin
              real_value= -6390;
              imag_value=32131;
            end
    10467 : begin
              real_value= -12784;
              imag_value=30163;
            end
    10468 : begin
              real_value= -18644;
              imag_value=26938;
            end
    10469 : begin
              real_value= -23726;
              imag_value=22589;
            end
    10470 : begin
              real_value= -27820;
              imag_value=17299;
            end
    10471 : begin
              real_value= -30755;
              imag_value=11289;
            end
    10472 : begin
              real_value= -32407;
              imag_value=4806;
            end
    10473 : begin
              real_value= -32707;
              imag_value=-1874;
            end
    10474 : begin
              real_value= -31645;
              imag_value=-8477;
            end
    10475 : begin
              real_value= -29263;
              imag_value=-14728;
            end
    10476 : begin
              real_value= -25661;
              imag_value=-20365;
            end
    10477 : begin
              real_value= -20988;
              imag_value=-25154;
            end
    10478 : begin
              real_value= -15442;
              imag_value=-28892;
            end
    10479 : begin
              real_value= -9253;
              imag_value=-31426;
            end
    10480 : begin
              real_value= -2676;
              imag_value=-32651;
            end
    10481 : begin
              real_value= 4009;
              imag_value=-32515;
            end
    10482 : begin
              real_value= 10529;
              imag_value=-31023;
            end
    10483 : begin
              real_value= 16611;
              imag_value=-28236;
            end
    10484 : begin
              real_value= 22001;
              imag_value=-24274;
            end
    10485 : begin
              real_value= 26472;
              imag_value=-19299;
            end
    10486 : begin
              real_value= 29841;
              imag_value=-13520;
            end
    10487 : begin
              real_value= 31965;
              imag_value=-7177;
            end
    10488 : begin
              real_value= 32757;
              imag_value=-535;
            end
    10489 : begin
              real_value= 32183;
              imag_value=6127;
            end
    10490 : begin
              real_value= 30267;
              imag_value=12537;
            end
    10491 : begin
              real_value= 27090;
              imag_value=18423;
            end
    10492 : begin
              real_value= 22782;
              imag_value=23541;
            end
    10493 : begin
              real_value= 17525;
              imag_value=27678;
            end
    10494 : begin
              real_value= 11539;
              imag_value=30661;
            end
    10495 : begin
              real_value= 5071;
              imag_value=32365;
            end
    10496 : begin
              real_value= -1606;
              imag_value=32721;
            end
    10497 : begin
              real_value= -8219;
              imag_value=31713;
            end
    10498 : begin
              real_value= -14489;
              imag_value=29382;
            end
    10499 : begin
              real_value= -20154;
              imag_value=25826;
            end
    10500 : begin
              real_value= -24981;
              imag_value=21194;
            end
    10501 : begin
              real_value= -28766;
              imag_value=15678;
            end
    10502 : begin
              real_value= -31351;
              imag_value=9508;
            end
    10503 : begin
              real_value= -32629;
              imag_value=2942;
            end
    10504 : begin
              real_value= -32547;
              imag_value=-3742;
            end
    10505 : begin
              real_value= -31107;
              imag_value=-10275;
            end
    10506 : begin
              real_value= -28371;
              imag_value=-16380;
            end
    10507 : begin
              real_value= -24453;
              imag_value=-21801;
            end
    10508 : begin
              real_value= -19515;
              imag_value=-26314;
            end
    10509 : begin
              real_value= -13764;
              imag_value=-29729;
            end
    10510 : begin
              real_value= -7438;
              imag_value=-31905;
            end
    10511 : begin
              real_value= -802;
              imag_value=-32750;
            end
    10512 : begin
              real_value= 5864;
              imag_value=-32231;
            end
    10513 : begin
              real_value= 12288;
              imag_value=-30369;
            end
    10514 : begin
              real_value= 18200;
              imag_value=-27240;
            end
    10515 : begin
              real_value= 23354;
              imag_value=-22974;
            end
    10516 : begin
              real_value= 27534;
              imag_value=-17752;
            end
    10517 : begin
              real_value= 30565;
              imag_value=-11790;
            end
    10518 : begin
              real_value= 32323;
              imag_value=-5336;
            end
    10519 : begin
              real_value= 32733;
              imag_value=1338;
            end
    10520 : begin
              real_value= 31779;
              imag_value=7959;
            end
    10521 : begin
              real_value= 29499;
              imag_value=14248;
            end
    10522 : begin
              real_value= 25990;
              imag_value=19943;
            end
    10523 : begin
              real_value= 21399;
              imag_value=24806;
            end
    10524 : begin
              real_value= 15914;
              imag_value=28636;
            end
    10525 : begin
              real_value= 9765;
              imag_value=31271;
            end
    10526 : begin
              real_value= 3210;
              imag_value=32603;
            end
    10527 : begin
              real_value= -3476;
              imag_value=32575;
            end
    10528 : begin
              real_value= -10021;
              imag_value=31191;
            end
    10529 : begin
              real_value= -16148;
              imag_value=28506;
            end
    10530 : begin
              real_value= -21600;
              imag_value=24630;
            end
    10531 : begin
              real_value= -26152;
              imag_value=19729;
            end
    10532 : begin
              real_value= -29615;
              imag_value=14006;
            end
    10533 : begin
              real_value= -31843;
              imag_value=7699;
            end
    10534 : begin
              real_value= -32743;
              imag_value=1070;
            end
    10535 : begin
              real_value= -32278;
              imag_value=-5599;
            end
    10536 : begin
              real_value= -30468;
              imag_value=-12039;
            end
    10537 : begin
              real_value= -27387;
              imag_value=-17977;
            end
    10538 : begin
              real_value= -23165;
              imag_value=-23165;
            end
    10539 : begin
              real_value= -17977;
              imag_value=-27387;
            end
    10540 : begin
              real_value= -12039;
              imag_value=-30468;
            end
    10541 : begin
              real_value= -5599;
              imag_value=-32278;
            end
    10542 : begin
              real_value= 1070;
              imag_value=-32743;
            end
    10543 : begin
              real_value= 7699;
              imag_value=-31843;
            end
    10544 : begin
              real_value= 14006;
              imag_value=-29615;
            end
    10545 : begin
              real_value= 19729;
              imag_value=-26152;
            end
    10546 : begin
              real_value= 24630;
              imag_value=-21600;
            end
    10547 : begin
              real_value= 28506;
              imag_value=-16148;
            end
    10548 : begin
              real_value= 31191;
              imag_value=-10021;
            end
    10549 : begin
              real_value= 32575;
              imag_value=-3476;
            end
    10550 : begin
              real_value= 32603;
              imag_value=3210;
            end
    10551 : begin
              real_value= 31271;
              imag_value=9765;
            end
    10552 : begin
              real_value= 28636;
              imag_value=15914;
            end
    10553 : begin
              real_value= 24806;
              imag_value=21399;
            end
    10554 : begin
              real_value= 19943;
              imag_value=25990;
            end
    10555 : begin
              real_value= 14248;
              imag_value=29499;
            end
    10556 : begin
              real_value= 7959;
              imag_value=31779;
            end
    10557 : begin
              real_value= 1338;
              imag_value=32733;
            end
    10558 : begin
              real_value= -5336;
              imag_value=32323;
            end
    10559 : begin
              real_value= -11790;
              imag_value=30565;
            end
    10560 : begin
              real_value= -17752;
              imag_value=27534;
            end
    10561 : begin
              real_value= -22974;
              imag_value=23354;
            end
    10562 : begin
              real_value= -27240;
              imag_value=18200;
            end
    10563 : begin
              real_value= -30369;
              imag_value=12288;
            end
    10564 : begin
              real_value= -32231;
              imag_value=5864;
            end
    10565 : begin
              real_value= -32750;
              imag_value=-802;
            end
    10566 : begin
              real_value= -31905;
              imag_value=-7438;
            end
    10567 : begin
              real_value= -29729;
              imag_value=-13764;
            end
    10568 : begin
              real_value= -26314;
              imag_value=-19515;
            end
    10569 : begin
              real_value= -21801;
              imag_value=-24453;
            end
    10570 : begin
              real_value= -16380;
              imag_value=-28371;
            end
    10571 : begin
              real_value= -10275;
              imag_value=-31107;
            end
    10572 : begin
              real_value= -3742;
              imag_value=-32547;
            end
    10573 : begin
              real_value= 2942;
              imag_value=-32629;
            end
    10574 : begin
              real_value= 9508;
              imag_value=-31351;
            end
    10575 : begin
              real_value= 15678;
              imag_value=-28766;
            end
    10576 : begin
              real_value= 21194;
              imag_value=-24981;
            end
    10577 : begin
              real_value= 25826;
              imag_value=-20154;
            end
    10578 : begin
              real_value= 29382;
              imag_value=-14489;
            end
    10579 : begin
              real_value= 31713;
              imag_value=-8219;
            end
    10580 : begin
              real_value= 32721;
              imag_value=-1606;
            end
    10581 : begin
              real_value= 32365;
              imag_value=5071;
            end
    10582 : begin
              real_value= 30661;
              imag_value=11539;
            end
    10583 : begin
              real_value= 27678;
              imag_value=17525;
            end
    10584 : begin
              real_value= 23541;
              imag_value=22782;
            end
    10585 : begin
              real_value= 18423;
              imag_value=27090;
            end
    10586 : begin
              real_value= 12537;
              imag_value=30267;
            end
    10587 : begin
              real_value= 6127;
              imag_value=32183;
            end
    10588 : begin
              real_value= -535;
              imag_value=32757;
            end
    10589 : begin
              real_value= -7177;
              imag_value=31965;
            end
    10590 : begin
              real_value= -13520;
              imag_value=29841;
            end
    10591 : begin
              real_value= -19299;
              imag_value=26472;
            end
    10592 : begin
              real_value= -24274;
              imag_value=22001;
            end
    10593 : begin
              real_value= -28236;
              imag_value=16611;
            end
    10594 : begin
              real_value= -31023;
              imag_value=10529;
            end
    10595 : begin
              real_value= -32515;
              imag_value=4009;
            end
    10596 : begin
              real_value= -32651;
              imag_value=-2676;
            end
    10597 : begin
              real_value= -31426;
              imag_value=-9253;
            end
    10598 : begin
              real_value= -28892;
              imag_value=-15442;
            end
    10599 : begin
              real_value= -25154;
              imag_value=-20988;
            end
    10600 : begin
              real_value= -20365;
              imag_value=-25661;
            end
    10601 : begin
              real_value= -14728;
              imag_value=-29263;
            end
    10602 : begin
              real_value= -8477;
              imag_value=-31645;
            end
    10603 : begin
              real_value= -1874;
              imag_value=-32707;
            end
    10604 : begin
              real_value= 4806;
              imag_value=-32407;
            end
    10605 : begin
              real_value= 11289;
              imag_value=-30755;
            end
    10606 : begin
              real_value= 17299;
              imag_value=-27820;
            end
    10607 : begin
              real_value= 22589;
              imag_value=-23726;
            end
    10608 : begin
              real_value= 26938;
              imag_value=-18644;
            end
    10609 : begin
              real_value= 30163;
              imag_value=-12784;
            end
    10610 : begin
              real_value= 32131;
              imag_value=-6390;
            end
    10611 : begin
              real_value= 32759;
              imag_value=267;
            end
    10612 : begin
              real_value= 32022;
              imag_value=6915;
            end
    10613 : begin
              real_value= 29950;
              imag_value=13274;
            end
    10614 : begin
              real_value= 26630;
              imag_value=19081;
            end
    10615 : begin
              real_value= 22199;
              imag_value=24092;
            end
    10616 : begin
              real_value= 16842;
              imag_value=28100;
            end
    10617 : begin
              real_value= 10783;
              imag_value=30935;
            end
    10618 : begin
              real_value= 4275;
              imag_value=32481;
            end
    10619 : begin
              real_value= -2408;
              imag_value=32673;
            end
    10620 : begin
              real_value= -8995;
              imag_value=31501;
            end
    10621 : begin
              real_value= -15206;
              imag_value=29017;
            end
    10622 : begin
              real_value= -20783;
              imag_value=25324;
            end
    10623 : begin
              real_value= -25494;
              imag_value=20575;
            end
    10624 : begin
              real_value= -29142;
              imag_value=14968;
            end
    10625 : begin
              real_value= -31575;
              imag_value=8737;
            end
    10626 : begin
              real_value= -32691;
              imag_value=2142;
            end
    10627 : begin
              real_value= -32445;
              imag_value=-4540;
            end
    10628 : begin
              real_value= -30846;
              imag_value=-11036;
            end
    10629 : begin
              real_value= -27961;
              imag_value=-17072;
            end
    10630 : begin
              real_value= -23911;
              imag_value=-22395;
            end
    10631 : begin
              real_value= -18863;
              imag_value=-26784;
            end
    10632 : begin
              real_value= -13030;
              imag_value=-30057;
            end
    10633 : begin
              real_value= -6654;
              imag_value=-32077;
            end
    10634 : begin
              real_value= 0;
              imag_value=-32760;
            end
    10635 : begin
              real_value= 6654;
              imag_value=-32077;
            end
    10636 : begin
              real_value= 13030;
              imag_value=-30057;
            end
    10637 : begin
              real_value= 18863;
              imag_value=-26784;
            end
    10638 : begin
              real_value= 23911;
              imag_value=-22395;
            end
    10639 : begin
              real_value= 27961;
              imag_value=-17072;
            end
    10640 : begin
              real_value= 30846;
              imag_value=-11036;
            end
    10641 : begin
              real_value= 32445;
              imag_value=-4540;
            end
    10642 : begin
              real_value= 32691;
              imag_value=2142;
            end
    10643 : begin
              real_value= 31575;
              imag_value=8737;
            end
    10644 : begin
              real_value= 29142;
              imag_value=14968;
            end
    10645 : begin
              real_value= 25494;
              imag_value=20575;
            end
    10646 : begin
              real_value= 20783;
              imag_value=25324;
            end
    10647 : begin
              real_value= 15206;
              imag_value=29017;
            end
    10648 : begin
              real_value= 8995;
              imag_value=31501;
            end
    10649 : begin
              real_value= 2408;
              imag_value=32673;
            end
    10650 : begin
              real_value= -4275;
              imag_value=32481;
            end
    10651 : begin
              real_value= -10783;
              imag_value=30935;
            end
    10652 : begin
              real_value= -16842;
              imag_value=28100;
            end
    10653 : begin
              real_value= -22199;
              imag_value=24092;
            end
    10654 : begin
              real_value= -26630;
              imag_value=19081;
            end
    10655 : begin
              real_value= -29950;
              imag_value=13274;
            end
    10656 : begin
              real_value= -32022;
              imag_value=6915;
            end
    10657 : begin
              real_value= -32759;
              imag_value=267;
            end
    10658 : begin
              real_value= -32131;
              imag_value=-6390;
            end
    10659 : begin
              real_value= -30163;
              imag_value=-12784;
            end
    10660 : begin
              real_value= -26938;
              imag_value=-18644;
            end
    10661 : begin
              real_value= -22589;
              imag_value=-23726;
            end
    10662 : begin
              real_value= -17299;
              imag_value=-27820;
            end
    10663 : begin
              real_value= -11289;
              imag_value=-30755;
            end
    10664 : begin
              real_value= -4806;
              imag_value=-32407;
            end
    10665 : begin
              real_value= 1874;
              imag_value=-32707;
            end
    10666 : begin
              real_value= 8477;
              imag_value=-31645;
            end
    10667 : begin
              real_value= 14728;
              imag_value=-29263;
            end
    10668 : begin
              real_value= 20365;
              imag_value=-25661;
            end
    10669 : begin
              real_value= 25154;
              imag_value=-20988;
            end
    10670 : begin
              real_value= 28892;
              imag_value=-15442;
            end
    10671 : begin
              real_value= 31426;
              imag_value=-9253;
            end
    10672 : begin
              real_value= 32651;
              imag_value=-2676;
            end
    10673 : begin
              real_value= 32515;
              imag_value=4009;
            end
    10674 : begin
              real_value= 31023;
              imag_value=10529;
            end
    10675 : begin
              real_value= 28236;
              imag_value=16611;
            end
    10676 : begin
              real_value= 24274;
              imag_value=22001;
            end
    10677 : begin
              real_value= 19299;
              imag_value=26472;
            end
    10678 : begin
              real_value= 13520;
              imag_value=29841;
            end
    10679 : begin
              real_value= 7177;
              imag_value=31965;
            end
    10680 : begin
              real_value= 535;
              imag_value=32757;
            end
    10681 : begin
              real_value= -6127;
              imag_value=32183;
            end
    10682 : begin
              real_value= -12537;
              imag_value=30267;
            end
    10683 : begin
              real_value= -18423;
              imag_value=27090;
            end
    10684 : begin
              real_value= -23541;
              imag_value=22782;
            end
    10685 : begin
              real_value= -27678;
              imag_value=17525;
            end
    10686 : begin
              real_value= -30661;
              imag_value=11539;
            end
    10687 : begin
              real_value= -32365;
              imag_value=5071;
            end
    10688 : begin
              real_value= -32721;
              imag_value=-1606;
            end
    10689 : begin
              real_value= -31713;
              imag_value=-8219;
            end
    10690 : begin
              real_value= -29382;
              imag_value=-14489;
            end
    10691 : begin
              real_value= -25826;
              imag_value=-20154;
            end
    10692 : begin
              real_value= -21194;
              imag_value=-24981;
            end
    10693 : begin
              real_value= -15678;
              imag_value=-28766;
            end
    10694 : begin
              real_value= -9508;
              imag_value=-31351;
            end
    10695 : begin
              real_value= -2942;
              imag_value=-32629;
            end
    10696 : begin
              real_value= 3742;
              imag_value=-32547;
            end
    10697 : begin
              real_value= 10275;
              imag_value=-31107;
            end
    10698 : begin
              real_value= 16380;
              imag_value=-28371;
            end
    10699 : begin
              real_value= 21801;
              imag_value=-24453;
            end
    10700 : begin
              real_value= 26314;
              imag_value=-19515;
            end
    10701 : begin
              real_value= 29729;
              imag_value=-13764;
            end
    10702 : begin
              real_value= 31905;
              imag_value=-7438;
            end
    10703 : begin
              real_value= 32750;
              imag_value=-802;
            end
    10704 : begin
              real_value= 32231;
              imag_value=5864;
            end
    10705 : begin
              real_value= 30369;
              imag_value=12288;
            end
    10706 : begin
              real_value= 27240;
              imag_value=18200;
            end
    10707 : begin
              real_value= 22974;
              imag_value=23354;
            end
    10708 : begin
              real_value= 17752;
              imag_value=27534;
            end
    10709 : begin
              real_value= 11790;
              imag_value=30565;
            end
    10710 : begin
              real_value= 5336;
              imag_value=32323;
            end
    10711 : begin
              real_value= -1338;
              imag_value=32733;
            end
    10712 : begin
              real_value= -7959;
              imag_value=31779;
            end
    10713 : begin
              real_value= -14248;
              imag_value=29499;
            end
    10714 : begin
              real_value= -19943;
              imag_value=25990;
            end
    10715 : begin
              real_value= -24806;
              imag_value=21399;
            end
    10716 : begin
              real_value= -28636;
              imag_value=15914;
            end
    10717 : begin
              real_value= -31271;
              imag_value=9765;
            end
    10718 : begin
              real_value= -32603;
              imag_value=3210;
            end
    10719 : begin
              real_value= -32575;
              imag_value=-3476;
            end
    10720 : begin
              real_value= -31191;
              imag_value=-10021;
            end
    10721 : begin
              real_value= -28506;
              imag_value=-16148;
            end
    10722 : begin
              real_value= -24630;
              imag_value=-21600;
            end
    10723 : begin
              real_value= -19729;
              imag_value=-26152;
            end
    10724 : begin
              real_value= -14006;
              imag_value=-29615;
            end
    10725 : begin
              real_value= -7699;
              imag_value=-31843;
            end
    10726 : begin
              real_value= -1070;
              imag_value=-32743;
            end
    10727 : begin
              real_value= 5599;
              imag_value=-32278;
            end
    10728 : begin
              real_value= 12039;
              imag_value=-30468;
            end
    10729 : begin
              real_value= 17977;
              imag_value=-27387;
            end
    10730 : begin
              real_value= 23165;
              imag_value=-23165;
            end
    10731 : begin
              real_value= 27387;
              imag_value=-17977;
            end
    10732 : begin
              real_value= 30468;
              imag_value=-12039;
            end
    10733 : begin
              real_value= 32278;
              imag_value=-5599;
            end
    10734 : begin
              real_value= 32743;
              imag_value=1070;
            end
    10735 : begin
              real_value= 31843;
              imag_value=7699;
            end
    10736 : begin
              real_value= 29615;
              imag_value=14006;
            end
    10737 : begin
              real_value= 26152;
              imag_value=19729;
            end
    10738 : begin
              real_value= 21600;
              imag_value=24630;
            end
    10739 : begin
              real_value= 16148;
              imag_value=28506;
            end
    10740 : begin
              real_value= 10021;
              imag_value=31191;
            end
    10741 : begin
              real_value= 3476;
              imag_value=32575;
            end
    10742 : begin
              real_value= -3210;
              imag_value=32603;
            end
    10743 : begin
              real_value= -9765;
              imag_value=31271;
            end
    10744 : begin
              real_value= -15914;
              imag_value=28636;
            end
    10745 : begin
              real_value= -21399;
              imag_value=24806;
            end
    10746 : begin
              real_value= -25990;
              imag_value=19943;
            end
    10747 : begin
              real_value= -29499;
              imag_value=14248;
            end
    10748 : begin
              real_value= -31779;
              imag_value=7959;
            end
    10749 : begin
              real_value= -32733;
              imag_value=1338;
            end
    10750 : begin
              real_value= -32323;
              imag_value=-5336;
            end
    10751 : begin
              real_value= -30565;
              imag_value=-11790;
            end
    10752 : begin
              real_value= -27534;
              imag_value=-17752;
            end
    10753 : begin
              real_value= -23354;
              imag_value=-22974;
            end
    10754 : begin
              real_value= -18200;
              imag_value=-27240;
            end
    10755 : begin
              real_value= -12288;
              imag_value=-30369;
            end
    10756 : begin
              real_value= -5864;
              imag_value=-32231;
            end
    10757 : begin
              real_value= 802;
              imag_value=-32750;
            end
    10758 : begin
              real_value= 7438;
              imag_value=-31905;
            end
    10759 : begin
              real_value= 13764;
              imag_value=-29729;
            end
    10760 : begin
              real_value= 19515;
              imag_value=-26314;
            end
    10761 : begin
              real_value= 24453;
              imag_value=-21801;
            end
    10762 : begin
              real_value= 28371;
              imag_value=-16380;
            end
    10763 : begin
              real_value= 31107;
              imag_value=-10275;
            end
    10764 : begin
              real_value= 32547;
              imag_value=-3742;
            end
    10765 : begin
              real_value= 32629;
              imag_value=2942;
            end
    10766 : begin
              real_value= 31351;
              imag_value=9508;
            end
    10767 : begin
              real_value= 28766;
              imag_value=15678;
            end
    10768 : begin
              real_value= 24981;
              imag_value=21194;
            end
    10769 : begin
              real_value= 20154;
              imag_value=25826;
            end
    10770 : begin
              real_value= 14489;
              imag_value=29382;
            end
    10771 : begin
              real_value= 8219;
              imag_value=31713;
            end
    10772 : begin
              real_value= 1606;
              imag_value=32721;
            end
    10773 : begin
              real_value= -5071;
              imag_value=32365;
            end
    10774 : begin
              real_value= -11539;
              imag_value=30661;
            end
    10775 : begin
              real_value= -17525;
              imag_value=27678;
            end
    10776 : begin
              real_value= -22782;
              imag_value=23541;
            end
    10777 : begin
              real_value= -27090;
              imag_value=18423;
            end
    10778 : begin
              real_value= -30267;
              imag_value=12537;
            end
    10779 : begin
              real_value= -32183;
              imag_value=6127;
            end
    10780 : begin
              real_value= -32757;
              imag_value=-535;
            end
    10781 : begin
              real_value= -31965;
              imag_value=-7177;
            end
    10782 : begin
              real_value= -29841;
              imag_value=-13520;
            end
    10783 : begin
              real_value= -26472;
              imag_value=-19299;
            end
    10784 : begin
              real_value= -22001;
              imag_value=-24274;
            end
    10785 : begin
              real_value= -16611;
              imag_value=-28236;
            end
    10786 : begin
              real_value= -10529;
              imag_value=-31023;
            end
    10787 : begin
              real_value= -4009;
              imag_value=-32515;
            end
    10788 : begin
              real_value= 2676;
              imag_value=-32651;
            end
    10789 : begin
              real_value= 9253;
              imag_value=-31426;
            end
    10790 : begin
              real_value= 15442;
              imag_value=-28892;
            end
    10791 : begin
              real_value= 20988;
              imag_value=-25154;
            end
    10792 : begin
              real_value= 25661;
              imag_value=-20365;
            end
    10793 : begin
              real_value= 29263;
              imag_value=-14728;
            end
    10794 : begin
              real_value= 31645;
              imag_value=-8477;
            end
    10795 : begin
              real_value= 32707;
              imag_value=-1874;
            end
    10796 : begin
              real_value= 32407;
              imag_value=4806;
            end
    10797 : begin
              real_value= 30755;
              imag_value=11289;
            end
    10798 : begin
              real_value= 27820;
              imag_value=17299;
            end
    10799 : begin
              real_value= 23726;
              imag_value=22589;
            end
    10800 : begin
              real_value= 18644;
              imag_value=26938;
            end
    10801 : begin
              real_value= 12784;
              imag_value=30163;
            end
    10802 : begin
              real_value= 6390;
              imag_value=32131;
            end
    10803 : begin
              real_value= -267;
              imag_value=32759;
            end
    10804 : begin
              real_value= -6915;
              imag_value=32022;
            end
    10805 : begin
              real_value= -13274;
              imag_value=29950;
            end
    10806 : begin
              real_value= -19081;
              imag_value=26630;
            end
    10807 : begin
              real_value= -24092;
              imag_value=22199;
            end
    10808 : begin
              real_value= -28100;
              imag_value=16842;
            end
    10809 : begin
              real_value= -30935;
              imag_value=10783;
            end
    10810 : begin
              real_value= -32481;
              imag_value=4275;
            end
    10811 : begin
              real_value= -32673;
              imag_value=-2408;
            end
    10812 : begin
              real_value= -31501;
              imag_value=-8995;
            end
    10813 : begin
              real_value= -29017;
              imag_value=-15206;
            end
    10814 : begin
              real_value= -25324;
              imag_value=-20783;
            end
    10815 : begin
              real_value= -20575;
              imag_value=-25494;
            end
    10816 : begin
              real_value= -14968;
              imag_value=-29142;
            end
    10817 : begin
              real_value= -8737;
              imag_value=-31575;
            end
    10818 : begin
              real_value= -2142;
              imag_value=-32691;
            end
    10819 : begin
              real_value= 4540;
              imag_value=-32445;
            end
    10820 : begin
              real_value= 11036;
              imag_value=-30846;
            end
    10821 : begin
              real_value= 17072;
              imag_value=-27961;
            end
    10822 : begin
              real_value= 22395;
              imag_value=-23911;
            end
    10823 : begin
              real_value= 26784;
              imag_value=-18863;
            end
    10824 : begin
              real_value= 30057;
              imag_value=-13030;
            end
    10825 : begin
              real_value= 32077;
              imag_value=-6654;
            end
    10826 : begin
              real_value= 32760;
              imag_value=0;
            end
    10827 : begin
              real_value= 32077;
              imag_value=6654;
            end
    10828 : begin
              real_value= 30057;
              imag_value=13030;
            end
    10829 : begin
              real_value= 26784;
              imag_value=18863;
            end
    10830 : begin
              real_value= 22395;
              imag_value=23911;
            end
    10831 : begin
              real_value= 17072;
              imag_value=27961;
            end
    10832 : begin
              real_value= 11036;
              imag_value=30846;
            end
    10833 : begin
              real_value= 4540;
              imag_value=32445;
            end
    10834 : begin
              real_value= -2142;
              imag_value=32691;
            end
    10835 : begin
              real_value= -8737;
              imag_value=31575;
            end
    10836 : begin
              real_value= -14968;
              imag_value=29142;
            end
    10837 : begin
              real_value= -20575;
              imag_value=25494;
            end
    10838 : begin
              real_value= -25324;
              imag_value=20783;
            end
    10839 : begin
              real_value= -29017;
              imag_value=15206;
            end
    10840 : begin
              real_value= -31501;
              imag_value=8995;
            end
    10841 : begin
              real_value= -32673;
              imag_value=2408;
            end
    10842 : begin
              real_value= -32481;
              imag_value=-4275;
            end
    10843 : begin
              real_value= -30935;
              imag_value=-10783;
            end
    10844 : begin
              real_value= -28100;
              imag_value=-16842;
            end
    10845 : begin
              real_value= -24092;
              imag_value=-22199;
            end
    10846 : begin
              real_value= -19081;
              imag_value=-26630;
            end
    10847 : begin
              real_value= -13274;
              imag_value=-29950;
            end
    10848 : begin
              real_value= -6915;
              imag_value=-32022;
            end
    10849 : begin
              real_value= -267;
              imag_value=-32759;
            end
    10850 : begin
              real_value= 6390;
              imag_value=-32131;
            end
    10851 : begin
              real_value= 12784;
              imag_value=-30163;
            end
    10852 : begin
              real_value= 18644;
              imag_value=-26938;
            end
    10853 : begin
              real_value= 23726;
              imag_value=-22589;
            end
    10854 : begin
              real_value= 27820;
              imag_value=-17299;
            end
    10855 : begin
              real_value= 30755;
              imag_value=-11289;
            end
    10856 : begin
              real_value= 32407;
              imag_value=-4806;
            end
    10857 : begin
              real_value= 32707;
              imag_value=1874;
            end
    10858 : begin
              real_value= 31645;
              imag_value=8477;
            end
    10859 : begin
              real_value= 29263;
              imag_value=14728;
            end
    10860 : begin
              real_value= 25661;
              imag_value=20365;
            end
    10861 : begin
              real_value= 20988;
              imag_value=25154;
            end
    10862 : begin
              real_value= 15442;
              imag_value=28892;
            end
    10863 : begin
              real_value= 9253;
              imag_value=31426;
            end
    10864 : begin
              real_value= 2676;
              imag_value=32651;
            end
    10865 : begin
              real_value= -4009;
              imag_value=32515;
            end
    10866 : begin
              real_value= -10529;
              imag_value=31023;
            end
    10867 : begin
              real_value= -16611;
              imag_value=28236;
            end
    10868 : begin
              real_value= -22001;
              imag_value=24274;
            end
    10869 : begin
              real_value= -26472;
              imag_value=19299;
            end
    10870 : begin
              real_value= -29841;
              imag_value=13520;
            end
    10871 : begin
              real_value= -31965;
              imag_value=7177;
            end
    10872 : begin
              real_value= -32757;
              imag_value=535;
            end
    10873 : begin
              real_value= -32183;
              imag_value=-6127;
            end
    10874 : begin
              real_value= -30267;
              imag_value=-12537;
            end
    10875 : begin
              real_value= -27090;
              imag_value=-18423;
            end
    10876 : begin
              real_value= -22782;
              imag_value=-23541;
            end
    10877 : begin
              real_value= -17525;
              imag_value=-27678;
            end
    10878 : begin
              real_value= -11539;
              imag_value=-30661;
            end
    10879 : begin
              real_value= -5071;
              imag_value=-32365;
            end
    10880 : begin
              real_value= 1606;
              imag_value=-32721;
            end
    10881 : begin
              real_value= 8219;
              imag_value=-31713;
            end
    10882 : begin
              real_value= 14489;
              imag_value=-29382;
            end
    10883 : begin
              real_value= 20154;
              imag_value=-25826;
            end
    10884 : begin
              real_value= 24981;
              imag_value=-21194;
            end
    10885 : begin
              real_value= 28766;
              imag_value=-15678;
            end
    10886 : begin
              real_value= 31351;
              imag_value=-9508;
            end
    10887 : begin
              real_value= 32629;
              imag_value=-2942;
            end
    10888 : begin
              real_value= 32547;
              imag_value=3742;
            end
    10889 : begin
              real_value= 31107;
              imag_value=10275;
            end
    10890 : begin
              real_value= 28371;
              imag_value=16380;
            end
    10891 : begin
              real_value= 24453;
              imag_value=21801;
            end
    10892 : begin
              real_value= 19515;
              imag_value=26314;
            end
    10893 : begin
              real_value= 13764;
              imag_value=29729;
            end
    10894 : begin
              real_value= 7438;
              imag_value=31905;
            end
    10895 : begin
              real_value= 802;
              imag_value=32750;
            end
    10896 : begin
              real_value= -5864;
              imag_value=32231;
            end
    10897 : begin
              real_value= -12288;
              imag_value=30369;
            end
    10898 : begin
              real_value= -18200;
              imag_value=27240;
            end
    10899 : begin
              real_value= -23354;
              imag_value=22974;
            end
    10900 : begin
              real_value= -27534;
              imag_value=17752;
            end
    10901 : begin
              real_value= -30565;
              imag_value=11790;
            end
    10902 : begin
              real_value= -32323;
              imag_value=5336;
            end
    10903 : begin
              real_value= -32733;
              imag_value=-1338;
            end
    10904 : begin
              real_value= -31779;
              imag_value=-7959;
            end
    10905 : begin
              real_value= -29499;
              imag_value=-14248;
            end
    10906 : begin
              real_value= -25990;
              imag_value=-19943;
            end
    10907 : begin
              real_value= -21399;
              imag_value=-24806;
            end
    10908 : begin
              real_value= -15914;
              imag_value=-28636;
            end
    10909 : begin
              real_value= -9765;
              imag_value=-31271;
            end
    10910 : begin
              real_value= -3210;
              imag_value=-32603;
            end
    10911 : begin
              real_value= 3476;
              imag_value=-32575;
            end
    10912 : begin
              real_value= 10021;
              imag_value=-31191;
            end
    10913 : begin
              real_value= 16148;
              imag_value=-28506;
            end
    10914 : begin
              real_value= 21600;
              imag_value=-24630;
            end
    10915 : begin
              real_value= 26152;
              imag_value=-19729;
            end
    10916 : begin
              real_value= 29615;
              imag_value=-14006;
            end
    10917 : begin
              real_value= 31843;
              imag_value=-7699;
            end
    10918 : begin
              real_value= 32743;
              imag_value=-1070;
            end
    10919 : begin
              real_value= 32278;
              imag_value=5599;
            end
    10920 : begin
              real_value= 30468;
              imag_value=12039;
            end
    10921 : begin
              real_value= 27387;
              imag_value=17977;
            end
    10922 : begin
              real_value= 23165;
              imag_value=23165;
            end
    10923 : begin
              real_value= 17977;
              imag_value=27387;
            end
    10924 : begin
              real_value= 12039;
              imag_value=30468;
            end
    10925 : begin
              real_value= 5599;
              imag_value=32278;
            end
    10926 : begin
              real_value= -1070;
              imag_value=32743;
            end
    10927 : begin
              real_value= -7699;
              imag_value=31843;
            end
    10928 : begin
              real_value= -14006;
              imag_value=29615;
            end
    10929 : begin
              real_value= -19729;
              imag_value=26152;
            end
    10930 : begin
              real_value= -24630;
              imag_value=21600;
            end
    10931 : begin
              real_value= -28506;
              imag_value=16148;
            end
    10932 : begin
              real_value= -31191;
              imag_value=10021;
            end
    10933 : begin
              real_value= -32575;
              imag_value=3476;
            end
    10934 : begin
              real_value= -32603;
              imag_value=-3210;
            end
    10935 : begin
              real_value= -31271;
              imag_value=-9765;
            end
    10936 : begin
              real_value= -28636;
              imag_value=-15914;
            end
    10937 : begin
              real_value= -24806;
              imag_value=-21399;
            end
    10938 : begin
              real_value= -19943;
              imag_value=-25990;
            end
    10939 : begin
              real_value= -14248;
              imag_value=-29499;
            end
    10940 : begin
              real_value= -7959;
              imag_value=-31779;
            end
    10941 : begin
              real_value= -1338;
              imag_value=-32733;
            end
    10942 : begin
              real_value= 5336;
              imag_value=-32323;
            end
    10943 : begin
              real_value= 11790;
              imag_value=-30565;
            end
    10944 : begin
              real_value= 17752;
              imag_value=-27534;
            end
    10945 : begin
              real_value= 22974;
              imag_value=-23354;
            end
    10946 : begin
              real_value= 27240;
              imag_value=-18200;
            end
    10947 : begin
              real_value= 30369;
              imag_value=-12288;
            end
    10948 : begin
              real_value= 32231;
              imag_value=-5864;
            end
    10949 : begin
              real_value= 32750;
              imag_value=802;
            end
    10950 : begin
              real_value= 31905;
              imag_value=7438;
            end
    10951 : begin
              real_value= 29729;
              imag_value=13764;
            end
    10952 : begin
              real_value= 26314;
              imag_value=19515;
            end
    10953 : begin
              real_value= 21801;
              imag_value=24453;
            end
    10954 : begin
              real_value= 16380;
              imag_value=28371;
            end
    10955 : begin
              real_value= 10275;
              imag_value=31107;
            end
    10956 : begin
              real_value= 3742;
              imag_value=32547;
            end
    10957 : begin
              real_value= -2942;
              imag_value=32629;
            end
    10958 : begin
              real_value= -9508;
              imag_value=31351;
            end
    10959 : begin
              real_value= -15678;
              imag_value=28766;
            end
    10960 : begin
              real_value= -21194;
              imag_value=24981;
            end
    10961 : begin
              real_value= -25826;
              imag_value=20154;
            end
    10962 : begin
              real_value= -29382;
              imag_value=14489;
            end
    10963 : begin
              real_value= -31713;
              imag_value=8219;
            end
    10964 : begin
              real_value= -32721;
              imag_value=1606;
            end
    10965 : begin
              real_value= -32365;
              imag_value=-5071;
            end
    10966 : begin
              real_value= -30661;
              imag_value=-11539;
            end
    10967 : begin
              real_value= -27678;
              imag_value=-17525;
            end
    10968 : begin
              real_value= -23541;
              imag_value=-22782;
            end
    10969 : begin
              real_value= -18423;
              imag_value=-27090;
            end
    10970 : begin
              real_value= -12537;
              imag_value=-30267;
            end
    10971 : begin
              real_value= -6127;
              imag_value=-32183;
            end
    10972 : begin
              real_value= 535;
              imag_value=-32757;
            end
    10973 : begin
              real_value= 7176;
              imag_value=-31965;
            end
    10974 : begin
              real_value= 13520;
              imag_value=-29841;
            end
    10975 : begin
              real_value= 19299;
              imag_value=-26473;
            end
    10976 : begin
              real_value= 24272;
              imag_value=-22000;
            end
    10977 : begin
              real_value= 28235;
              imag_value=-16611;
            end
    10978 : begin
              real_value= 31023;
              imag_value=-10531;
            end
    10979 : begin
              real_value= 32513;
              imag_value=-4009;
            end
    10980 : begin
              real_value= 32649;
              imag_value=2676;
            end
    10981 : begin
              real_value= 31429;
              imag_value=9250;
            end
    10982 : begin
              real_value= 28893;
              imag_value=15441;
            end
    10983 : begin
              real_value= 25149;
              imag_value=20990;
            end
    10984 : begin
              real_value= 20369;
              imag_value=25658;
            end
    10985 : begin
              real_value= 14732;
              imag_value=29261;
            end
    10986 : begin
              real_value= 8470;
              imag_value=31649;
            end
    10987 : begin
              real_value= 1874;
              imag_value=32706;
            end
    10988 : begin
              real_value= -4796;
              imag_value=32401;
            end
    10989 : begin
              real_value= -11296;
              imag_value=30760;
            end
    10990 : begin
              real_value= -17306;
              imag_value=27822;
            end
    10991 : begin
              real_value= -22575;
              imag_value=23717;
            end
    10992 : begin
              real_value= -26942;
              imag_value=18647;
            end
    10993 : begin
              real_value= -30180;
              imag_value=12791;
            end
    10994 : begin
              real_value= -32115;
              imag_value=6379;
            end
    10995 : begin
              real_value= -32752;
              imag_value=-270;
            end
    10996 : begin
              real_value= -32048;
              imag_value=-6901;
            end
    10997 : begin
              real_value= -29939;
              imag_value=-13284;
            end
    10998 : begin
              real_value= -26606;
              imag_value=-19093;
            end
    10999 : begin
              real_value= -22231;
              imag_value=-24074;
            end
    11000 : begin
              real_value= -16848;
              imag_value=-28101;
            end
    11001 : begin
              real_value= -10741;
              imag_value=-30958;
            end
    11002 : begin
              real_value= -4302;
              imag_value=-32463;
            end
    11003 : begin
              real_value= 2376;
              imag_value=-32659;
            end
    11004 : begin
              real_value= 9050;
              imag_value=-31535;
            end
    11005 : begin
              real_value= 15203;
              imag_value=-29011;
            end
    11006 : begin
              real_value= 20718;
              imag_value=-25291;
            end
    11007 : begin
              real_value= 25545;
              imag_value=-20610;
            end
    11008 : begin
              real_value= 29180;
              imag_value=-14983;
            end
    11009 : begin
              real_value= 31485;
              imag_value=-8686;
            end
    11010 : begin
              real_value= 32713;
              imag_value=-2164;
            end
    11011 : begin
              real_value= 32536;
              imag_value=4494;
            end
    11012 : begin
              real_value= 30753;
              imag_value=11095;
            end
    11013 : begin
              real_value= 27924;
              imag_value=17081;
            end
    11014 : begin
              real_value= 24049;
              imag_value=22318;
            end
    11015 : begin
              real_value= 18805;
              imag_value=26830;
            end
    11016 : begin
              real_value= 12912;
              imag_value=30113;
            end
    11017 : begin
              real_value= 6813;
              imag_value=31982;
            end
    11018 : begin
              real_value= 22;
              imag_value=32766;
            end
    11019 : begin
              real_value= -6857;
              imag_value=32187;
            end
    11020 : begin
              real_value= -12904;
              imag_value=29970;
            end
    11021 : begin
              real_value= -18716;
              imag_value=26721;
            end
    11022 : begin
              real_value= -24171;
              imag_value=22548;
            end
    11023 : begin
              real_value= -27943;
              imag_value=17034;
            end
    11024 : begin
              real_value= -30550;
              imag_value=10883;
            end
    11025 : begin
              real_value= -32693;
              imag_value=4703;
            end
    11026 : begin
              real_value= -32767;
              imag_value=-2079;
            end
    11027 : begin
              real_value= -31143;
              imag_value=-8983;
            end
    11028 : begin
              real_value= -29265;
              imag_value=-14857;
            end
    11029 : begin
              real_value= -25945;
              imag_value=-20355;
            end
    11030 : begin
              real_value= -20279;
              imag_value=-25639;
            end
    11031 : begin
              real_value= -15027;
              imag_value=-29056;
            end
    11032 : begin
              real_value= -9820;
              imag_value=-31056;
            end
    11033 : begin
              real_value= -1975;
              imag_value=-32767;
            end
    11034 : begin
              real_value= 5098;
              imag_value=-32767;
            end
    11035 : begin
              real_value= 9346;
              imag_value=-30107;
            end
    11036 : begin
              real_value= 16836;
              imag_value=-28276;
            end
    11037 : begin
              real_value= 25291;
              imag_value=-25624;
            end
    11038 : begin
              real_value= 21019;
              imag_value=-15986;
            end
    11039 : begin
              real_value= 5512;
              imag_value=-3264;
            end
    11040 : begin
              real_value= -2886;
              imag_value=1887;
            end
    11041 : begin
              real_value= -148;
              imag_value=-93;
            end
    11042 : begin
              real_value= 1441;
              imag_value=-817;
            end
    11043 : begin
              real_value= -738;
              imag_value=518;
            end
    11044 : begin
              real_value= -495;
              imag_value=209;
            end
    11045 : begin
              real_value= 801;
              imag_value=-484;
            end
    11046 : begin
              real_value= -122;
              imag_value=134;
            end
    11047 : begin
              real_value= -526;
              imag_value=273;
            end
    11048 : begin
              real_value= 417;
              imag_value=-276;
            end
    11049 : begin
              real_value= 157;
              imag_value=-48;
            end
    11050 : begin
              real_value= -429;
              imag_value=246;
            end
    11051 : begin
              real_value= 142;
              imag_value=-116;
            end
    11052 : begin
              real_value= 265;
              imag_value=-130;
            end
    11053 : begin
              real_value= -280;
              imag_value=176;
            end
    11054 : begin
              real_value= -40;
              imag_value=-2;
            end
    11055 : begin
              real_value= 263;
              imag_value=-145;
            end
    11056 : begin
              real_value= -128;
              imag_value=94;
            end
    11057 : begin
              real_value= -138;
              imag_value=63;
            end
    11058 : begin
              real_value= 196;
              imag_value=-118;
            end
    11059 : begin
              real_value= -5;
              imag_value=22;
            end
    11060 : begin
              real_value= -162;
              imag_value=87;
            end
    11061 : begin
              real_value= 107;
              imag_value=-72;
            end
    11062 : begin
              real_value= 67;
              imag_value=-25;
            end
    11063 : begin
              real_value= -135;
              imag_value=79;
            end
    11064 : begin
              real_value= 25;
              imag_value=-25;
            end
    11065 : begin
              real_value= 96;
              imag_value=-49;
            end
    11066 : begin
              real_value= -84;
              imag_value=54;
            end
    11067 : begin
              real_value= -29;
              imag_value=6;
            end
    11068 : begin
              real_value= 88;
              imag_value=-50;
            end
    11069 : begin
              real_value= -31;
              imag_value=24;
            end
    11070 : begin
              real_value= -55;
              imag_value=25;
            end
    11071 : begin
              real_value= 60;
              imag_value=-38;
            end
    11072 : begin
              real_value= 6;
              imag_value=0;
            end
    11073 : begin
              real_value= -55;
              imag_value=29;
            end
    11074 : begin
              real_value= 26;
              imag_value=-20;
            end
    11075 : begin
              real_value= 27;
              imag_value=-12;
            end
    11076 : begin
              real_value= -40;
              imag_value=23;
            end
    11077 : begin
              real_value= 1;
              imag_value=-4;
            end
    11078 : begin
              real_value= 31;
              imag_value=-17;
            end
    11079 : begin
              real_value= -20;
              imag_value=13;
            end
    11080 : begin
              real_value= -12;
              imag_value=3;
            end
    11081 : begin
              real_value= 24;
              imag_value=-14;
            end
    11082 : begin
              real_value= -4;
              imag_value=3;
            end
    11083 : begin
              real_value= -16;
              imag_value=7;
            end
    11084 : begin
              real_value= 13;
              imag_value=-9;
            end
    11085 : begin
              real_value= 3;
              imag_value=0;
            end
    11086 : begin
              real_value= -13;
              imag_value=6;
            end
    11087 : begin
              real_value= 4;
              imag_value=-3;
            end
    11088 : begin
              real_value= 7;
              imag_value=-3;
            end
    11089 : begin
              real_value= -8;
              imag_value=4;
            end
    11090 : begin
              real_value= 0;
              imag_value=0;
            end
    11091 : begin
              real_value= 6;
              imag_value=-3;
            end
    11092 : begin
              real_value= -2;
              imag_value=1;
            end
    11093 : begin
              real_value= -3;
              imag_value=0;
            end
    11094 : begin
              real_value= 2;
              imag_value=-2;
            end
    11095 : begin
              real_value= 0;
              imag_value=0;
            end
    11096 : begin
              real_value= -2;
              imag_value=0;
            end
    11097 : begin
              real_value= 0;
              imag_value=-1;
            end
    11098 : begin
              real_value= 0;
              imag_value=0;
            end
    11099 : begin
              real_value= 0;
              imag_value=0;
            end
    11100 : begin
              real_value= 0;
              imag_value=0;
            end
    11101 : begin
              real_value= 0;
              imag_value=0;
            end
    11102 : begin
              real_value= 0;
              imag_value=0;
            end
    11103 : begin
              real_value= 0;
              imag_value=0;
            end
    11104 : begin
              real_value= 0;
              imag_value=0;
            end
    11105 : begin
              real_value= 0;
              imag_value=0;
            end
    11106 : begin
              real_value= 0;
              imag_value=0;
            end
    11107 : begin
              real_value= 0;
              imag_value=0;
            end
    11108 : begin
              real_value= 0;
              imag_value=0;
            end
    11109 : begin
              real_value= 0;
              imag_value=0;
            end
    11110 : begin
              real_value= 0;
              imag_value=0;
            end
    11111 : begin
              real_value= 0;
              imag_value=0;
            end
    11112 : begin
              real_value= 0;
              imag_value=0;
            end
    11113 : begin
              real_value= 0;
              imag_value=0;
            end
    11114 : begin
              real_value= 0;
              imag_value=0;
            end
    11115 : begin
              real_value= 0;
              imag_value=0;
            end
    11116 : begin
              real_value= 0;
              imag_value=0;
            end
    11117 : begin
              real_value= 0;
              imag_value=0;
            end
    11118 : begin
              real_value= 0;
              imag_value=0;
            end
    11119 : begin
              real_value= 0;
              imag_value=0;
            end
    11120 : begin
              real_value= 0;
              imag_value=0;
            end
    11121 : begin
              real_value= 0;
              imag_value=0;
            end
    11122 : begin
              real_value= 0;
              imag_value=0;
            end
    11123 : begin
              real_value= 0;
              imag_value=0;
            end
    11124 : begin
              real_value= 0;
              imag_value=0;
            end
    11125 : begin
              real_value= 0;
              imag_value=0;
            end
    11126 : begin
              real_value= 0;
              imag_value=0;
            end
    11127 : begin
              real_value= 0;
              imag_value=0;
            end
    11128 : begin
              real_value= 0;
              imag_value=0;
            end
    11129 : begin
              real_value= 0;
              imag_value=0;
            end
    11130 : begin
              real_value= 0;
              imag_value=0;
            end
    11131 : begin
              real_value= 0;
              imag_value=0;
            end
    11132 : begin
              real_value= 0;
              imag_value=0;
            end
    11133 : begin
              real_value= 0;
              imag_value=0;
            end
    11134 : begin
              real_value= 0;
              imag_value=0;
            end
    11135 : begin
              real_value= 0;
              imag_value=0;
            end
    11136 : begin
              real_value= 0;
              imag_value=0;
            end
    11137 : begin
              real_value= 0;
              imag_value=0;
            end
    11138 : begin
              real_value= 0;
              imag_value=0;
            end
    11139 : begin
              real_value= 0;
              imag_value=0;
            end
    11140 : begin
              real_value= 0;
              imag_value=0;
            end
    11141 : begin
              real_value= 0;
              imag_value=0;
            end
    11142 : begin
              real_value= 0;
              imag_value=0;
            end
    11143 : begin
              real_value= 0;
              imag_value=0;
            end
    11144 : begin
              real_value= 0;
              imag_value=0;
            end
    11145 : begin
              real_value= 0;
              imag_value=0;
            end
    11146 : begin
              real_value= 0;
              imag_value=0;
            end
    11147 : begin
              real_value= 0;
              imag_value=0;
            end
    11148 : begin
              real_value= 0;
              imag_value=0;
            end
    11149 : begin
              real_value= 0;
              imag_value=0;
            end
    11150 : begin
              real_value= 0;
              imag_value=0;
            end
    11151 : begin
              real_value= 0;
              imag_value=0;
            end
    11152 : begin
              real_value= 0;
              imag_value=0;
            end
    11153 : begin
              real_value= 0;
              imag_value=0;
            end
    11154 : begin
              real_value= 0;
              imag_value=0;
            end
    11155 : begin
              real_value= 0;
              imag_value=0;
            end
    11156 : begin
              real_value= 0;
              imag_value=0;
            end
    11157 : begin
              real_value= 0;
              imag_value=0;
            end
    11158 : begin
              real_value= 0;
              imag_value=0;
            end
    11159 : begin
              real_value= 0;
              imag_value=0;
            end
    11160 : begin
              real_value= 0;
              imag_value=0;
            end
    11161 : begin
              real_value= 0;
              imag_value=0;
            end
    11162 : begin
              real_value= 0;
              imag_value=0;
            end
    11163 : begin
              real_value= 0;
              imag_value=0;
            end
    11164 : begin
              real_value= 0;
              imag_value=0;
            end
    11165 : begin
              real_value= 0;
              imag_value=0;
            end
    11166 : begin
              real_value= 0;
              imag_value=0;
            end
    11167 : begin
              real_value= 0;
              imag_value=0;
            end
    11168 : begin
              real_value= 0;
              imag_value=0;
            end
    11169 : begin
              real_value= 0;
              imag_value=0;
            end
    11170 : begin
              real_value= 0;
              imag_value=0;
            end
    11171 : begin
              real_value= 0;
              imag_value=0;
            end
    11172 : begin
              real_value= 0;
              imag_value=0;
            end
    11173 : begin
              real_value= 0;
              imag_value=0;
            end
    11174 : begin
              real_value= 0;
              imag_value=0;
            end
    11175 : begin
              real_value= 0;
              imag_value=0;
            end
    11176 : begin
              real_value= 0;
              imag_value=0;
            end
    11177 : begin
              real_value= 0;
              imag_value=0;
            end
    11178 : begin
              real_value= 0;
              imag_value=0;
            end
    11179 : begin
              real_value= 0;
              imag_value=0;
            end
    11180 : begin
              real_value= 0;
              imag_value=0;
            end
    11181 : begin
              real_value= 0;
              imag_value=0;
            end
    11182 : begin
              real_value= 0;
              imag_value=0;
            end
    11183 : begin
              real_value= 0;
              imag_value=0;
            end
    11184 : begin
              real_value= 0;
              imag_value=0;
            end
    11185 : begin
              real_value= 0;
              imag_value=0;
            end
    11186 : begin
              real_value= 0;
              imag_value=0;
            end
    11187 : begin
              real_value= 0;
              imag_value=0;
            end
    11188 : begin
              real_value= 0;
              imag_value=0;
            end
    11189 : begin
              real_value= 0;
              imag_value=0;
            end
    11190 : begin
              real_value= 0;
              imag_value=0;
            end
    11191 : begin
              real_value= 0;
              imag_value=0;
            end
    11192 : begin
              real_value= 0;
              imag_value=0;
            end
    11193 : begin
              real_value= 0;
              imag_value=0;
            end
    11194 : begin
              real_value= 0;
              imag_value=0;
            end
    11195 : begin
              real_value= 0;
              imag_value=0;
            end
    11196 : begin
              real_value= 0;
              imag_value=0;
            end
    11197 : begin
              real_value= 0;
              imag_value=0;
            end
    11198 : begin
              real_value= 0;
              imag_value=0;
            end
    11199 : begin
              real_value= 0;
              imag_value=0;
            end
    11200 : begin
              real_value= 0;
              imag_value=0;
            end
    11201 : begin
              real_value= 0;
              imag_value=0;
            end
    11202 : begin
              real_value= 0;
              imag_value=0;
            end
    11203 : begin
              real_value= 0;
              imag_value=0;
            end
    11204 : begin
              real_value= 0;
              imag_value=0;
            end
    11205 : begin
              real_value= 0;
              imag_value=0;
            end
    11206 : begin
              real_value= 0;
              imag_value=0;
            end
    11207 : begin
              real_value= 0;
              imag_value=0;
            end
    11208 : begin
              real_value= 0;
              imag_value=0;
            end
    11209 : begin
              real_value= 0;
              imag_value=0;
            end
    11210 : begin
              real_value= 0;
              imag_value=0;
            end
    11211 : begin
              real_value= 0;
              imag_value=0;
            end
    11212 : begin
              real_value= 0;
              imag_value=0;
            end
    11213 : begin
              real_value= 0;
              imag_value=0;
            end
    11214 : begin
              real_value= 0;
              imag_value=0;
            end
    11215 : begin
              real_value= 0;
              imag_value=0;
            end
    11216 : begin
              real_value= 0;
              imag_value=0;
            end
    11217 : begin
              real_value= 0;
              imag_value=0;
            end
    11218 : begin
              real_value= 0;
              imag_value=0;
            end
    11219 : begin
              real_value= 0;
              imag_value=0;
            end
    11220 : begin
              real_value= 0;
              imag_value=0;
            end
    11221 : begin
              real_value= 0;
              imag_value=0;
            end
    11222 : begin
              real_value= 0;
              imag_value=0;
            end
    11223 : begin
              real_value= 0;
              imag_value=0;
            end
    11224 : begin
              real_value= 0;
              imag_value=0;
            end
    11225 : begin
              real_value= 0;
              imag_value=0;
            end
    11226 : begin
              real_value= 0;
              imag_value=0;
            end
    11227 : begin
              real_value= 0;
              imag_value=0;
            end
    11228 : begin
              real_value= 0;
              imag_value=0;
            end
    11229 : begin
              real_value= 0;
              imag_value=0;
            end
    11230 : begin
              real_value= 0;
              imag_value=0;
            end
    11231 : begin
              real_value= 0;
              imag_value=0;
            end
    11232 : begin
              real_value= 0;
              imag_value=0;
            end
    11233 : begin
              real_value= 0;
              imag_value=0;
            end
    11234 : begin
              real_value= 0;
              imag_value=0;
            end
    11235 : begin
              real_value= 0;
              imag_value=0;
            end
    11236 : begin
              real_value= 0;
              imag_value=0;
            end
    11237 : begin
              real_value= 0;
              imag_value=0;
            end
    11238 : begin
              real_value= 0;
              imag_value=0;
            end
    11239 : begin
              real_value= 0;
              imag_value=0;
            end
    11240 : begin
              real_value= 0;
              imag_value=0;
            end
    11241 : begin
              real_value= 0;
              imag_value=0;
            end
    11242 : begin
              real_value= 0;
              imag_value=0;
            end
    11243 : begin
              real_value= 0;
              imag_value=0;
            end
    11244 : begin
              real_value= 0;
              imag_value=0;
            end
    11245 : begin
              real_value= 0;
              imag_value=0;
            end
    11246 : begin
              real_value= 0;
              imag_value=0;
            end
    11247 : begin
              real_value= 0;
              imag_value=0;
            end
    11248 : begin
              real_value= 0;
              imag_value=0;
            end
    11249 : begin
              real_value= 0;
              imag_value=0;
            end
    11250 : begin
              real_value= 0;
              imag_value=0;
            end
    11251 : begin
              real_value= 0;
              imag_value=0;
            end
    11252 : begin
              real_value= 0;
              imag_value=0;
            end
    11253 : begin
              real_value= 0;
              imag_value=0;
            end
    11254 : begin
              real_value= 0;
              imag_value=0;
            end
    11255 : begin
              real_value= 0;
              imag_value=0;
            end
    11256 : begin
              real_value= 0;
              imag_value=0;
            end
    11257 : begin
              real_value= 0;
              imag_value=0;
            end
    11258 : begin
              real_value= 0;
              imag_value=0;
            end
    11259 : begin
              real_value= 0;
              imag_value=0;
            end
    11260 : begin
              real_value= 0;
              imag_value=0;
            end
    11261 : begin
              real_value= 0;
              imag_value=0;
            end
    11262 : begin
              real_value= 0;
              imag_value=0;
            end
    11263 : begin
              real_value= 0;
              imag_value=0;
            end
    11264 : begin
              real_value= 0;
              imag_value=0;
            end
    11265 : begin
              real_value= 0;
              imag_value=0;
            end
    11266 : begin
              real_value= 0;
              imag_value=0;
            end
    11267 : begin
              real_value= 0;
              imag_value=0;
            end
    11268 : begin
              real_value= 0;
              imag_value=0;
            end
    11269 : begin
              real_value= 0;
              imag_value=0;
            end
    11270 : begin
              real_value= 0;
              imag_value=0;
            end
    11271 : begin
              real_value= 0;
              imag_value=0;
            end
    11272 : begin
              real_value= 0;
              imag_value=0;
            end
    11273 : begin
              real_value= 0;
              imag_value=0;
            end
    11274 : begin
              real_value= 0;
              imag_value=0;
            end
    11275 : begin
              real_value= 0;
              imag_value=0;
            end
    11276 : begin
              real_value= 0;
              imag_value=0;
            end
    11277 : begin
              real_value= 0;
              imag_value=0;
            end
    11278 : begin
              real_value= 0;
              imag_value=0;
            end
    11279 : begin
              real_value= 0;
              imag_value=0;
            end
    11280 : begin
              real_value= 0;
              imag_value=0;
            end
    11281 : begin
              real_value= 0;
              imag_value=0;
            end
    11282 : begin
              real_value= 0;
              imag_value=0;
            end
    11283 : begin
              real_value= 0;
              imag_value=0;
            end
    11284 : begin
              real_value= 0;
              imag_value=0;
            end
    11285 : begin
              real_value= 0;
              imag_value=0;
            end
    11286 : begin
              real_value= 0;
              imag_value=0;
            end
    11287 : begin
              real_value= 0;
              imag_value=0;
            end
    11288 : begin
              real_value= 0;
              imag_value=0;
            end
    11289 : begin
              real_value= 0;
              imag_value=0;
            end
    11290 : begin
              real_value= 0;
              imag_value=0;
            end
    11291 : begin
              real_value= 0;
              imag_value=0;
            end
    11292 : begin
              real_value= 0;
              imag_value=0;
            end
    11293 : begin
              real_value= 0;
              imag_value=0;
            end
    11294 : begin
              real_value= 0;
              imag_value=0;
            end
    11295 : begin
              real_value= 0;
              imag_value=0;
            end
    11296 : begin
              real_value= 0;
              imag_value=0;
            end
    11297 : begin
              real_value= 0;
              imag_value=0;
            end
    11298 : begin
              real_value= 0;
              imag_value=0;
            end
    11299 : begin
              real_value= 0;
              imag_value=0;
            end
    11300 : begin
              real_value= 0;
              imag_value=0;
            end
    11301 : begin
              real_value= 0;
              imag_value=0;
            end
    11302 : begin
              real_value= 0;
              imag_value=0;
            end
    11303 : begin
              real_value= 0;
              imag_value=0;
            end
    11304 : begin
              real_value= 0;
              imag_value=0;
            end
    11305 : begin
              real_value= 0;
              imag_value=0;
            end
    11306 : begin
              real_value= 0;
              imag_value=0;
            end
    11307 : begin
              real_value= 0;
              imag_value=0;
            end
    11308 : begin
              real_value= 0;
              imag_value=0;
            end
    11309 : begin
              real_value= 0;
              imag_value=0;
            end
    11310 : begin
              real_value= 0;
              imag_value=0;
            end
    11311 : begin
              real_value= 0;
              imag_value=0;
            end
    11312 : begin
              real_value= 0;
              imag_value=0;
            end
    11313 : begin
              real_value= 0;
              imag_value=0;
            end
    11314 : begin
              real_value= 0;
              imag_value=0;
            end
    11315 : begin
              real_value= 0;
              imag_value=0;
            end
    11316 : begin
              real_value= 0;
              imag_value=0;
            end
    11317 : begin
              real_value= 0;
              imag_value=0;
            end
    11318 : begin
              real_value= 0;
              imag_value=0;
            end
    11319 : begin
              real_value= 0;
              imag_value=0;
            end
    11320 : begin
              real_value= 0;
              imag_value=0;
            end
    11321 : begin
              real_value= 0;
              imag_value=0;
            end
    11322 : begin
              real_value= 0;
              imag_value=0;
            end
    11323 : begin
              real_value= 0;
              imag_value=0;
            end
    11324 : begin
              real_value= 0;
              imag_value=0;
            end
    11325 : begin
              real_value= 0;
              imag_value=0;
            end
    11326 : begin
              real_value= 0;
              imag_value=0;
            end
    11327 : begin
              real_value= 0;
              imag_value=0;
            end
    11328 : begin
              real_value= 0;
              imag_value=0;
            end
    11329 : begin
              real_value= 0;
              imag_value=0;
            end
    11330 : begin
              real_value= 0;
              imag_value=0;
            end
    11331 : begin
              real_value= 0;
              imag_value=0;
            end
    11332 : begin
              real_value= 0;
              imag_value=0;
            end
    11333 : begin
              real_value= 0;
              imag_value=0;
            end
    11334 : begin
              real_value= 0;
              imag_value=0;
            end
    11335 : begin
              real_value= 0;
              imag_value=0;
            end
    11336 : begin
              real_value= 0;
              imag_value=0;
            end
    11337 : begin
              real_value= 0;
              imag_value=0;
            end
    11338 : begin
              real_value= 0;
              imag_value=0;
            end
    11339 : begin
              real_value= 0;
              imag_value=0;
            end
    11340 : begin
              real_value= 0;
              imag_value=0;
            end
    11341 : begin
              real_value= 0;
              imag_value=0;
            end
    11342 : begin
              real_value= 0;
              imag_value=0;
            end
    11343 : begin
              real_value= 0;
              imag_value=0;
            end
    11344 : begin
              real_value= 0;
              imag_value=0;
            end
    11345 : begin
              real_value= 0;
              imag_value=0;
            end
    11346 : begin
              real_value= 0;
              imag_value=0;
            end
    11347 : begin
              real_value= 0;
              imag_value=0;
            end
    11348 : begin
              real_value= 0;
              imag_value=0;
            end
    11349 : begin
              real_value= 0;
              imag_value=0;
            end
    11350 : begin
              real_value= 0;
              imag_value=0;
            end
    11351 : begin
              real_value= 0;
              imag_value=0;
            end
    11352 : begin
              real_value= 0;
              imag_value=0;
            end
    11353 : begin
              real_value= 0;
              imag_value=0;
            end
    11354 : begin
              real_value= 0;
              imag_value=0;
            end
    11355 : begin
              real_value= 0;
              imag_value=0;
            end
    11356 : begin
              real_value= 0;
              imag_value=0;
            end
    11357 : begin
              real_value= 0;
              imag_value=0;
            end
    11358 : begin
              real_value= 0;
              imag_value=0;
            end
    11359 : begin
              real_value= 0;
              imag_value=0;
            end
    11360 : begin
              real_value= 0;
              imag_value=0;
            end
    11361 : begin
              real_value= 0;
              imag_value=0;
            end
    11362 : begin
              real_value= 0;
              imag_value=0;
            end
    11363 : begin
              real_value= 0;
              imag_value=0;
            end
    11364 : begin
              real_value= 0;
              imag_value=0;
            end
    11365 : begin
              real_value= 0;
              imag_value=0;
            end
    11366 : begin
              real_value= 0;
              imag_value=0;
            end
    11367 : begin
              real_value= 0;
              imag_value=0;
            end
    11368 : begin
              real_value= 0;
              imag_value=0;
            end
    11369 : begin
              real_value= 0;
              imag_value=0;
            end
    11370 : begin
              real_value= 0;
              imag_value=0;
            end
    11371 : begin
              real_value= 0;
              imag_value=0;
            end
    11372 : begin
              real_value= 0;
              imag_value=0;
            end
    11373 : begin
              real_value= 0;
              imag_value=0;
            end
    11374 : begin
              real_value= 0;
              imag_value=0;
            end
    11375 : begin
              real_value= 0;
              imag_value=0;
            end
    11376 : begin
              real_value= 0;
              imag_value=0;
            end
    11377 : begin
              real_value= 0;
              imag_value=0;
            end
    11378 : begin
              real_value= 0;
              imag_value=0;
            end
    11379 : begin
              real_value= 0;
              imag_value=0;
            end
    11380 : begin
              real_value= 0;
              imag_value=0;
            end
    11381 : begin
              real_value= 0;
              imag_value=0;
            end
    11382 : begin
              real_value= 0;
              imag_value=0;
            end
    11383 : begin
              real_value= 0;
              imag_value=0;
            end
    11384 : begin
              real_value= 0;
              imag_value=0;
            end
    11385 : begin
              real_value= 0;
              imag_value=0;
            end
    11386 : begin
              real_value= 0;
              imag_value=0;
            end
    11387 : begin
              real_value= 0;
              imag_value=0;
            end
    11388 : begin
              real_value= 0;
              imag_value=0;
            end
    11389 : begin
              real_value= 0;
              imag_value=0;
            end
    11390 : begin
              real_value= 0;
              imag_value=0;
            end
    11391 : begin
              real_value= 0;
              imag_value=0;
            end
    11392 : begin
              real_value= 0;
              imag_value=0;
            end
    11393 : begin
              real_value= 0;
              imag_value=0;
            end
    11394 : begin
              real_value= 0;
              imag_value=0;
            end
    11395 : begin
              real_value= 0;
              imag_value=0;
            end
    11396 : begin
              real_value= 0;
              imag_value=0;
            end
    11397 : begin
              real_value= 0;
              imag_value=0;
            end
    11398 : begin
              real_value= 0;
              imag_value=0;
            end
    11399 : begin
              real_value= 0;
              imag_value=0;
            end
    11400 : begin
              real_value= 0;
              imag_value=0;
            end
    11401 : begin
              real_value= 0;
              imag_value=0;
            end
    11402 : begin
              real_value= 0;
              imag_value=0;
            end
    11403 : begin
              real_value= 0;
              imag_value=0;
            end
    11404 : begin
              real_value= 0;
              imag_value=0;
            end
    11405 : begin
              real_value= 0;
              imag_value=0;
            end
    11406 : begin
              real_value= 0;
              imag_value=0;
            end
    11407 : begin
              real_value= 0;
              imag_value=0;
            end
    11408 : begin
              real_value= 0;
              imag_value=0;
            end
    11409 : begin
              real_value= 0;
              imag_value=0;
            end
    11410 : begin
              real_value= 0;
              imag_value=0;
            end
    11411 : begin
              real_value= 0;
              imag_value=0;
            end
    11412 : begin
              real_value= 0;
              imag_value=0;
            end
    11413 : begin
              real_value= 0;
              imag_value=0;
            end
    11414 : begin
              real_value= 0;
              imag_value=0;
            end
    11415 : begin
              real_value= 0;
              imag_value=0;
            end
    11416 : begin
              real_value= 0;
              imag_value=0;
            end
    11417 : begin
              real_value= 0;
              imag_value=0;
            end
    11418 : begin
              real_value= 0;
              imag_value=0;
            end
    11419 : begin
              real_value= 0;
              imag_value=0;
            end
    11420 : begin
              real_value= 0;
              imag_value=0;
            end
    11421 : begin
              real_value= 0;
              imag_value=0;
            end
    11422 : begin
              real_value= 0;
              imag_value=0;
            end
    11423 : begin
              real_value= 0;
              imag_value=0;
            end
    11424 : begin
              real_value= 0;
              imag_value=0;
            end
    11425 : begin
              real_value= 0;
              imag_value=0;
            end
    11426 : begin
              real_value= 0;
              imag_value=0;
            end
    11427 : begin
              real_value= 0;
              imag_value=0;
            end
    11428 : begin
              real_value= 0;
              imag_value=0;
            end
    11429 : begin
              real_value= 0;
              imag_value=0;
            end
    11430 : begin
              real_value= 0;
              imag_value=0;
            end
    11431 : begin
              real_value= 0;
              imag_value=0;
            end
    11432 : begin
              real_value= 0;
              imag_value=0;
            end
    11433 : begin
              real_value= 0;
              imag_value=0;
            end
    11434 : begin
              real_value= 0;
              imag_value=0;
            end
    11435 : begin
              real_value= 0;
              imag_value=0;
            end
    11436 : begin
              real_value= 0;
              imag_value=0;
            end
    11437 : begin
              real_value= 0;
              imag_value=0;
            end
    11438 : begin
              real_value= 0;
              imag_value=0;
            end
    11439 : begin
              real_value= 0;
              imag_value=0;
            end
    11440 : begin
              real_value= 0;
              imag_value=0;
            end
    11441 : begin
              real_value= 0;
              imag_value=0;
            end
    11442 : begin
              real_value= 0;
              imag_value=0;
            end
    11443 : begin
              real_value= 0;
              imag_value=0;
            end
    11444 : begin
              real_value= 0;
              imag_value=0;
            end
    11445 : begin
              real_value= 0;
              imag_value=0;
            end
    11446 : begin
              real_value= 0;
              imag_value=0;
            end
    11447 : begin
              real_value= 0;
              imag_value=0;
            end
    11448 : begin
              real_value= 0;
              imag_value=0;
            end
    11449 : begin
              real_value= 0;
              imag_value=0;
            end
    11450 : begin
              real_value= 0;
              imag_value=0;
            end
    11451 : begin
              real_value= 0;
              imag_value=0;
            end
    11452 : begin
              real_value= 0;
              imag_value=0;
            end
    11453 : begin
              real_value= 0;
              imag_value=0;
            end
    11454 : begin
              real_value= 0;
              imag_value=0;
            end
    11455 : begin
              real_value= 0;
              imag_value=0;
            end
    11456 : begin
              real_value= 0;
              imag_value=0;
            end
    11457 : begin
              real_value= 0;
              imag_value=0;
            end
    11458 : begin
              real_value= 0;
              imag_value=0;
            end
    11459 : begin
              real_value= 0;
              imag_value=0;
            end
    11460 : begin
              real_value= 0;
              imag_value=0;
            end
    11461 : begin
              real_value= 0;
              imag_value=0;
            end
    11462 : begin
              real_value= 0;
              imag_value=0;
            end
    11463 : begin
              real_value= 0;
              imag_value=0;
            end
    11464 : begin
              real_value= 0;
              imag_value=0;
            end
    11465 : begin
              real_value= 0;
              imag_value=0;
            end
    11466 : begin
              real_value= 0;
              imag_value=0;
            end
    11467 : begin
              real_value= 0;
              imag_value=0;
            end
    11468 : begin
              real_value= 0;
              imag_value=0;
            end
    11469 : begin
              real_value= 0;
              imag_value=0;
            end
    11470 : begin
              real_value= 0;
              imag_value=0;
            end
    11471 : begin
              real_value= 0;
              imag_value=0;
            end
    11472 : begin
              real_value= 0;
              imag_value=0;
            end
    11473 : begin
              real_value= 0;
              imag_value=0;
            end
    11474 : begin
              real_value= 0;
              imag_value=0;
            end
    11475 : begin
              real_value= 0;
              imag_value=0;
            end
    11476 : begin
              real_value= 0;
              imag_value=0;
            end
    11477 : begin
              real_value= 0;
              imag_value=0;
            end
    11478 : begin
              real_value= 0;
              imag_value=0;
            end
    11479 : begin
              real_value= 0;
              imag_value=0;
            end
    11480 : begin
              real_value= 0;
              imag_value=0;
            end
    11481 : begin
              real_value= 0;
              imag_value=0;
            end
    11482 : begin
              real_value= 0;
              imag_value=0;
            end
    11483 : begin
              real_value= 0;
              imag_value=0;
            end
    11484 : begin
              real_value= 0;
              imag_value=0;
            end
    11485 : begin
              real_value= 0;
              imag_value=0;
            end
    11486 : begin
              real_value= 0;
              imag_value=0;
            end
    11487 : begin
              real_value= 0;
              imag_value=0;
            end
    11488 : begin
              real_value= 0;
              imag_value=0;
            end
    11489 : begin
              real_value= 0;
              imag_value=0;
            end
    11490 : begin
              real_value= 0;
              imag_value=0;
            end
    11491 : begin
              real_value= 0;
              imag_value=0;
            end
    11492 : begin
              real_value= 0;
              imag_value=0;
            end
    11493 : begin
              real_value= 0;
              imag_value=0;
            end
    11494 : begin
              real_value= 0;
              imag_value=0;
            end
    11495 : begin
              real_value= 0;
              imag_value=0;
            end
    11496 : begin
              real_value= 0;
              imag_value=0;
            end
    11497 : begin
              real_value= 0;
              imag_value=0;
            end
    11498 : begin
              real_value= 0;
              imag_value=0;
            end
    11499 : begin
              real_value= 0;
              imag_value=0;
            end
    11500 : begin
              real_value= 0;
              imag_value=0;
            end
    11501 : begin
              real_value= 0;
              imag_value=0;
            end
    11502 : begin
              real_value= 0;
              imag_value=0;
            end
    11503 : begin
              real_value= 0;
              imag_value=0;
            end
    11504 : begin
              real_value= 0;
              imag_value=0;
            end
    11505 : begin
              real_value= 0;
              imag_value=0;
            end
    11506 : begin
              real_value= 0;
              imag_value=0;
            end
    11507 : begin
              real_value= 0;
              imag_value=0;
            end
    11508 : begin
              real_value= 0;
              imag_value=0;
            end
    11509 : begin
              real_value= 0;
              imag_value=0;
            end
    11510 : begin
              real_value= 0;
              imag_value=0;
            end
    11511 : begin
              real_value= 0;
              imag_value=0;
            end
    11512 : begin
              real_value= 0;
              imag_value=0;
            end
    11513 : begin
              real_value= 0;
              imag_value=0;
            end
    11514 : begin
              real_value= 0;
              imag_value=0;
            end
    11515 : begin
              real_value= 0;
              imag_value=0;
            end
    11516 : begin
              real_value= 0;
              imag_value=0;
            end
    11517 : begin
              real_value= 0;
              imag_value=0;
            end
    11518 : begin
              real_value= 0;
              imag_value=0;
            end
    11519 : begin
              real_value= 0;
              imag_value=0;
            end
    11520 : begin
              real_value= 0;
              imag_value=0;
            end
    11521 : begin
              real_value= 0;
              imag_value=0;
            end
    11522 : begin
              real_value= 0;
              imag_value=0;
            end
    11523 : begin
              real_value= 0;
              imag_value=0;
            end
    11524 : begin
              real_value= 0;
              imag_value=0;
            end
    11525 : begin
              real_value= 0;
              imag_value=0;
            end
    11526 : begin
              real_value= 0;
              imag_value=0;
            end
    11527 : begin
              real_value= 0;
              imag_value=0;
            end
    11528 : begin
              real_value= 0;
              imag_value=0;
            end
    11529 : begin
              real_value= 0;
              imag_value=0;
            end
    11530 : begin
              real_value= 0;
              imag_value=0;
            end
    11531 : begin
              real_value= 0;
              imag_value=0;
            end
    11532 : begin
              real_value= 0;
              imag_value=0;
            end
    11533 : begin
              real_value= 0;
              imag_value=0;
            end
    11534 : begin
              real_value= 0;
              imag_value=0;
            end
    11535 : begin
              real_value= 0;
              imag_value=0;
            end
    11536 : begin
              real_value= 0;
              imag_value=0;
            end
    11537 : begin
              real_value= 0;
              imag_value=0;
            end
    11538 : begin
              real_value= 0;
              imag_value=0;
            end
    11539 : begin
              real_value= 0;
              imag_value=0;
            end
    11540 : begin
              real_value= 0;
              imag_value=0;
            end
    11541 : begin
              real_value= 0;
              imag_value=0;
            end
    11542 : begin
              real_value= 0;
              imag_value=0;
            end
    11543 : begin
              real_value= 0;
              imag_value=0;
            end
    11544 : begin
              real_value= 0;
              imag_value=0;
            end
    11545 : begin
              real_value= 0;
              imag_value=0;
            end
    11546 : begin
              real_value= 0;
              imag_value=0;
            end
    11547 : begin
              real_value= 0;
              imag_value=0;
            end
    11548 : begin
              real_value= 0;
              imag_value=0;
            end
    11549 : begin
              real_value= 0;
              imag_value=0;
            end
    11550 : begin
              real_value= 0;
              imag_value=0;
            end
    11551 : begin
              real_value= 0;
              imag_value=0;
            end
    11552 : begin
              real_value= 0;
              imag_value=0;
            end
    11553 : begin
              real_value= 0;
              imag_value=0;
            end
    11554 : begin
              real_value= 0;
              imag_value=0;
            end
    11555 : begin
              real_value= 0;
              imag_value=0;
            end
    11556 : begin
              real_value= 0;
              imag_value=0;
            end
    11557 : begin
              real_value= 0;
              imag_value=0;
            end
    11558 : begin
              real_value= 0;
              imag_value=0;
            end
    11559 : begin
              real_value= 0;
              imag_value=0;
            end
    11560 : begin
              real_value= 0;
              imag_value=0;
            end
    11561 : begin
              real_value= 0;
              imag_value=0;
            end
    11562 : begin
              real_value= 0;
              imag_value=0;
            end
    11563 : begin
              real_value= 0;
              imag_value=0;
            end
    11564 : begin
              real_value= 0;
              imag_value=0;
            end
    11565 : begin
              real_value= 0;
              imag_value=0;
            end
    11566 : begin
              real_value= 0;
              imag_value=0;
            end
    11567 : begin
              real_value= 0;
              imag_value=0;
            end
    11568 : begin
              real_value= 0;
              imag_value=0;
            end
    11569 : begin
              real_value= 0;
              imag_value=0;
            end
    11570 : begin
              real_value= 0;
              imag_value=0;
            end
    11571 : begin
              real_value= 0;
              imag_value=0;
            end
    11572 : begin
              real_value= 0;
              imag_value=0;
            end
    11573 : begin
              real_value= 0;
              imag_value=0;
            end
    11574 : begin
              real_value= 0;
              imag_value=0;
            end
    11575 : begin
              real_value= 0;
              imag_value=0;
            end
    11576 : begin
              real_value= 0;
              imag_value=0;
            end
    11577 : begin
              real_value= 0;
              imag_value=0;
            end
    11578 : begin
              real_value= 0;
              imag_value=0;
            end
    11579 : begin
              real_value= 0;
              imag_value=0;
            end
    11580 : begin
              real_value= 0;
              imag_value=0;
            end
    11581 : begin
              real_value= 0;
              imag_value=0;
            end
    11582 : begin
              real_value= 0;
              imag_value=0;
            end
    11583 : begin
              real_value= 0;
              imag_value=0;
            end
    11584 : begin
              real_value= 0;
              imag_value=0;
            end
    11585 : begin
              real_value= 0;
              imag_value=0;
            end
    11586 : begin
              real_value= 0;
              imag_value=0;
            end
    11587 : begin
              real_value= 0;
              imag_value=0;
            end
    11588 : begin
              real_value= 0;
              imag_value=0;
            end
    11589 : begin
              real_value= 0;
              imag_value=0;
            end
    11590 : begin
              real_value= 0;
              imag_value=0;
            end
    11591 : begin
              real_value= 0;
              imag_value=0;
            end
    11592 : begin
              real_value= 0;
              imag_value=0;
            end
    11593 : begin
              real_value= 0;
              imag_value=0;
            end
    11594 : begin
              real_value= 0;
              imag_value=0;
            end
    11595 : begin
              real_value= 0;
              imag_value=0;
            end
    11596 : begin
              real_value= 0;
              imag_value=0;
            end
    11597 : begin
              real_value= 0;
              imag_value=0;
            end
    11598 : begin
              real_value= 0;
              imag_value=0;
            end
    11599 : begin
              real_value= 0;
              imag_value=0;
            end
    11600 : begin
              real_value= 0;
              imag_value=0;
            end
    11601 : begin
              real_value= 0;
              imag_value=0;
            end
    11602 : begin
              real_value= 0;
              imag_value=0;
            end
    11603 : begin
              real_value= 0;
              imag_value=0;
            end
    11604 : begin
              real_value= 0;
              imag_value=0;
            end
    11605 : begin
              real_value= 0;
              imag_value=0;
            end
    11606 : begin
              real_value= 0;
              imag_value=0;
            end
    11607 : begin
              real_value= 0;
              imag_value=0;
            end
    11608 : begin
              real_value= 0;
              imag_value=0;
            end
    11609 : begin
              real_value= 0;
              imag_value=0;
            end
    11610 : begin
              real_value= 0;
              imag_value=0;
            end
    11611 : begin
              real_value= 0;
              imag_value=0;
            end
    11612 : begin
              real_value= 0;
              imag_value=0;
            end
    11613 : begin
              real_value= 0;
              imag_value=0;
            end
    11614 : begin
              real_value= 0;
              imag_value=0;
            end
    11615 : begin
              real_value= 0;
              imag_value=0;
            end
    11616 : begin
              real_value= 0;
              imag_value=0;
            end
    11617 : begin
              real_value= 0;
              imag_value=0;
            end
    11618 : begin
              real_value= 0;
              imag_value=0;
            end
    11619 : begin
              real_value= 0;
              imag_value=0;
            end
    11620 : begin
              real_value= 0;
              imag_value=0;
            end
    11621 : begin
              real_value= 0;
              imag_value=0;
            end
    11622 : begin
              real_value= 0;
              imag_value=0;
            end
    11623 : begin
              real_value= 0;
              imag_value=0;
            end
    11624 : begin
              real_value= 0;
              imag_value=0;
            end
    11625 : begin
              real_value= 0;
              imag_value=0;
            end
    11626 : begin
              real_value= 0;
              imag_value=0;
            end
    11627 : begin
              real_value= 0;
              imag_value=0;
            end
    11628 : begin
              real_value= 0;
              imag_value=0;
            end
    11629 : begin
              real_value= 0;
              imag_value=0;
            end
    11630 : begin
              real_value= 0;
              imag_value=0;
            end
    11631 : begin
              real_value= 0;
              imag_value=0;
            end
    11632 : begin
              real_value= 0;
              imag_value=0;
            end
    11633 : begin
              real_value= 0;
              imag_value=0;
            end
    11634 : begin
              real_value= 0;
              imag_value=0;
            end
    11635 : begin
              real_value= 0;
              imag_value=0;
            end
    11636 : begin
              real_value= 0;
              imag_value=0;
            end
    11637 : begin
              real_value= 0;
              imag_value=0;
            end
    11638 : begin
              real_value= 0;
              imag_value=0;
            end
    11639 : begin
              real_value= 0;
              imag_value=0;
            end
    11640 : begin
              real_value= 0;
              imag_value=0;
            end
    11641 : begin
              real_value= 0;
              imag_value=0;
            end
    11642 : begin
              real_value= 0;
              imag_value=0;
            end
    11643 : begin
              real_value= 0;
              imag_value=0;
            end
    11644 : begin
              real_value= 0;
              imag_value=0;
            end
    11645 : begin
              real_value= 0;
              imag_value=0;
            end
    11646 : begin
              real_value= 0;
              imag_value=0;
            end
    11647 : begin
              real_value= 0;
              imag_value=0;
            end
    11648 : begin
              real_value= 0;
              imag_value=0;
            end
    11649 : begin
              real_value= 0;
              imag_value=0;
            end
    11650 : begin
              real_value= 0;
              imag_value=0;
            end
    11651 : begin
              real_value= 0;
              imag_value=0;
            end
    11652 : begin
              real_value= 0;
              imag_value=0;
            end
    11653 : begin
              real_value= 0;
              imag_value=0;
            end
    11654 : begin
              real_value= 0;
              imag_value=0;
            end
    11655 : begin
              real_value= 0;
              imag_value=0;
            end
    11656 : begin
              real_value= 0;
              imag_value=0;
            end
    11657 : begin
              real_value= 0;
              imag_value=0;
            end
    11658 : begin
              real_value= 0;
              imag_value=0;
            end
    11659 : begin
              real_value= 0;
              imag_value=0;
            end
    11660 : begin
              real_value= 0;
              imag_value=0;
            end
    11661 : begin
              real_value= 0;
              imag_value=0;
            end
    11662 : begin
              real_value= 0;
              imag_value=0;
            end
    11663 : begin
              real_value= 0;
              imag_value=0;
            end
    11664 : begin
              real_value= 0;
              imag_value=0;
            end
    11665 : begin
              real_value= 0;
              imag_value=0;
            end
    11666 : begin
              real_value= 0;
              imag_value=0;
            end
    11667 : begin
              real_value= 0;
              imag_value=0;
            end
    11668 : begin
              real_value= 0;
              imag_value=0;
            end
    11669 : begin
              real_value= 0;
              imag_value=0;
            end
    11670 : begin
              real_value= 0;
              imag_value=0;
            end
    11671 : begin
              real_value= 0;
              imag_value=0;
            end
    11672 : begin
              real_value= 0;
              imag_value=0;
            end
    11673 : begin
              real_value= 0;
              imag_value=0;
            end
    11674 : begin
              real_value= 0;
              imag_value=0;
            end
    11675 : begin
              real_value= 0;
              imag_value=0;
            end
    11676 : begin
              real_value= 0;
              imag_value=0;
            end
    11677 : begin
              real_value= 0;
              imag_value=0;
            end
    11678 : begin
              real_value= 0;
              imag_value=0;
            end
    11679 : begin
              real_value= 0;
              imag_value=0;
            end
    11680 : begin
              real_value= 0;
              imag_value=0;
            end
    11681 : begin
              real_value= 0;
              imag_value=0;
            end
    11682 : begin
              real_value= 0;
              imag_value=0;
            end
    11683 : begin
              real_value= 0;
              imag_value=0;
            end
    11684 : begin
              real_value= 0;
              imag_value=0;
            end
    11685 : begin
              real_value= 0;
              imag_value=0;
            end
    11686 : begin
              real_value= 0;
              imag_value=0;
            end
    11687 : begin
              real_value= 0;
              imag_value=0;
            end
    11688 : begin
              real_value= 0;
              imag_value=0;
            end
    11689 : begin
              real_value= 0;
              imag_value=0;
            end
    11690 : begin
              real_value= 0;
              imag_value=0;
            end
    11691 : begin
              real_value= 0;
              imag_value=0;
            end
    11692 : begin
              real_value= 0;
              imag_value=0;
            end
    11693 : begin
              real_value= 0;
              imag_value=0;
            end
    11694 : begin
              real_value= 0;
              imag_value=0;
            end
    11695 : begin
              real_value= 0;
              imag_value=0;
            end
    11696 : begin
              real_value= 0;
              imag_value=0;
            end
    11697 : begin
              real_value= 0;
              imag_value=0;
            end
    11698 : begin
              real_value= 0;
              imag_value=0;
            end
    11699 : begin
              real_value= 0;
              imag_value=0;
            end
    11700 : begin
              real_value= 0;
              imag_value=0;
            end
    11701 : begin
              real_value= 0;
              imag_value=0;
            end
    11702 : begin
              real_value= 0;
              imag_value=0;
            end
    11703 : begin
              real_value= 0;
              imag_value=0;
            end
    11704 : begin
              real_value= 0;
              imag_value=0;
            end
    11705 : begin
              real_value= 0;
              imag_value=0;
            end
    11706 : begin
              real_value= 0;
              imag_value=0;
            end
    11707 : begin
              real_value= 0;
              imag_value=0;
            end
    11708 : begin
              real_value= 0;
              imag_value=0;
            end
    11709 : begin
              real_value= 0;
              imag_value=0;
            end
    11710 : begin
              real_value= 0;
              imag_value=0;
            end
    11711 : begin
              real_value= 0;
              imag_value=0;
            end
    11712 : begin
              real_value= 0;
              imag_value=0;
            end
    11713 : begin
              real_value= 0;
              imag_value=0;
            end
    11714 : begin
              real_value= 0;
              imag_value=0;
            end
    11715 : begin
              real_value= 0;
              imag_value=0;
            end
    11716 : begin
              real_value= 0;
              imag_value=0;
            end
    11717 : begin
              real_value= 0;
              imag_value=0;
            end
    11718 : begin
              real_value= 0;
              imag_value=0;
            end
    11719 : begin
              real_value= 0;
              imag_value=0;
            end
    11720 : begin
              real_value= 0;
              imag_value=0;
            end
    11721 : begin
              real_value= 0;
              imag_value=0;
            end
    11722 : begin
              real_value= 0;
              imag_value=0;
            end
    11723 : begin
              real_value= 0;
              imag_value=0;
            end
    11724 : begin
              real_value= 0;
              imag_value=0;
            end
    11725 : begin
              real_value= 0;
              imag_value=0;
            end
    11726 : begin
              real_value= 0;
              imag_value=0;
            end
    11727 : begin
              real_value= 0;
              imag_value=0;
            end
    11728 : begin
              real_value= 0;
              imag_value=0;
            end
    11729 : begin
              real_value= 0;
              imag_value=0;
            end
    11730 : begin
              real_value= 0;
              imag_value=0;
            end
    11731 : begin
              real_value= 0;
              imag_value=0;
            end
    11732 : begin
              real_value= 0;
              imag_value=0;
            end
    11733 : begin
              real_value= 0;
              imag_value=0;
            end
    11734 : begin
              real_value= 0;
              imag_value=0;
            end
    11735 : begin
              real_value= 0;
              imag_value=0;
            end
    11736 : begin
              real_value= 0;
              imag_value=0;
            end
    11737 : begin
              real_value= 0;
              imag_value=0;
            end
    11738 : begin
              real_value= 0;
              imag_value=0;
            end
    11739 : begin
              real_value= 0;
              imag_value=0;
            end
    11740 : begin
              real_value= 0;
              imag_value=0;
            end
    11741 : begin
              real_value= 0;
              imag_value=0;
            end
    11742 : begin
              real_value= 0;
              imag_value=0;
            end
    11743 : begin
              real_value= 0;
              imag_value=0;
            end
    11744 : begin
              real_value= 0;
              imag_value=0;
            end
    11745 : begin
              real_value= 0;
              imag_value=0;
            end
    11746 : begin
              real_value= 0;
              imag_value=0;
            end
    11747 : begin
              real_value= 0;
              imag_value=0;
            end
    11748 : begin
              real_value= 0;
              imag_value=0;
            end
    11749 : begin
              real_value= 0;
              imag_value=0;
            end
    11750 : begin
              real_value= 0;
              imag_value=0;
            end
    11751 : begin
              real_value= 0;
              imag_value=0;
            end
    11752 : begin
              real_value= 0;
              imag_value=0;
            end
    11753 : begin
              real_value= 0;
              imag_value=0;
            end
    11754 : begin
              real_value= 0;
              imag_value=0;
            end
    11755 : begin
              real_value= 0;
              imag_value=0;
            end
    11756 : begin
              real_value= 0;
              imag_value=0;
            end
    11757 : begin
              real_value= 0;
              imag_value=0;
            end
    11758 : begin
              real_value= 0;
              imag_value=0;
            end
    11759 : begin
              real_value= 0;
              imag_value=0;
            end
    11760 : begin
              real_value= 0;
              imag_value=0;
            end
    11761 : begin
              real_value= 0;
              imag_value=0;
            end
    11762 : begin
              real_value= 0;
              imag_value=0;
            end
    11763 : begin
              real_value= 0;
              imag_value=0;
            end
    11764 : begin
              real_value= 0;
              imag_value=0;
            end
    11765 : begin
              real_value= 0;
              imag_value=0;
            end
    11766 : begin
              real_value= 0;
              imag_value=0;
            end
    11767 : begin
              real_value= 0;
              imag_value=0;
            end
    11768 : begin
              real_value= 0;
              imag_value=0;
            end
    11769 : begin
              real_value= 0;
              imag_value=0;
            end
    11770 : begin
              real_value= 0;
              imag_value=0;
            end
    11771 : begin
              real_value= 0;
              imag_value=0;
            end
    11772 : begin
              real_value= 0;
              imag_value=0;
            end
    11773 : begin
              real_value= 0;
              imag_value=0;
            end
    11774 : begin
              real_value= 0;
              imag_value=0;
            end
    11775 : begin
              real_value= 0;
              imag_value=0;
            end
    11776 : begin
              real_value= 0;
              imag_value=0;
            end
    11777 : begin
              real_value= 0;
              imag_value=0;
            end
    11778 : begin
              real_value= 0;
              imag_value=0;
            end
    11779 : begin
              real_value= 0;
              imag_value=0;
            end
    11780 : begin
              real_value= 0;
              imag_value=0;
            end
    11781 : begin
              real_value= 0;
              imag_value=0;
            end
    11782 : begin
              real_value= 0;
              imag_value=0;
            end
    11783 : begin
              real_value= 0;
              imag_value=0;
            end
    11784 : begin
              real_value= 0;
              imag_value=0;
            end
    11785 : begin
              real_value= 0;
              imag_value=0;
            end
    11786 : begin
              real_value= 0;
              imag_value=0;
            end
    11787 : begin
              real_value= 0;
              imag_value=0;
            end
    11788 : begin
              real_value= 0;
              imag_value=0;
            end
    11789 : begin
              real_value= 0;
              imag_value=0;
            end
    11790 : begin
              real_value= 0;
              imag_value=0;
            end
    11791 : begin
              real_value= 0;
              imag_value=0;
            end
    11792 : begin
              real_value= 0;
              imag_value=0;
            end
    11793 : begin
              real_value= 0;
              imag_value=0;
            end
    11794 : begin
              real_value= 0;
              imag_value=0;
            end
    11795 : begin
              real_value= 0;
              imag_value=0;
            end
    11796 : begin
              real_value= 0;
              imag_value=0;
            end
    11797 : begin
              real_value= 0;
              imag_value=0;
            end
    11798 : begin
              real_value= 0;
              imag_value=0;
            end
    11799 : begin
              real_value= 0;
              imag_value=0;
            end
    11800 : begin
              real_value= 0;
              imag_value=0;
            end
    11801 : begin
              real_value= 0;
              imag_value=0;
            end
    11802 : begin
              real_value= 0;
              imag_value=0;
            end
    11803 : begin
              real_value= 0;
              imag_value=0;
            end
    11804 : begin
              real_value= 0;
              imag_value=0;
            end
    11805 : begin
              real_value= 0;
              imag_value=0;
            end
    11806 : begin
              real_value= 0;
              imag_value=0;
            end
    11807 : begin
              real_value= 0;
              imag_value=0;
            end
    11808 : begin
              real_value= 0;
              imag_value=0;
            end
    11809 : begin
              real_value= 0;
              imag_value=0;
            end
    11810 : begin
              real_value= 0;
              imag_value=0;
            end
    11811 : begin
              real_value= 0;
              imag_value=0;
            end
    11812 : begin
              real_value= 0;
              imag_value=0;
            end
    11813 : begin
              real_value= 0;
              imag_value=0;
            end
    11814 : begin
              real_value= 0;
              imag_value=0;
            end
    11815 : begin
              real_value= 0;
              imag_value=0;
            end
    11816 : begin
              real_value= 0;
              imag_value=0;
            end
    11817 : begin
              real_value= 0;
              imag_value=0;
            end
    11818 : begin
              real_value= 0;
              imag_value=0;
            end
    11819 : begin
              real_value= 0;
              imag_value=0;
            end
    11820 : begin
              real_value= 0;
              imag_value=0;
            end
    11821 : begin
              real_value= 0;
              imag_value=0;
            end
    11822 : begin
              real_value= 0;
              imag_value=0;
            end
    11823 : begin
              real_value= 0;
              imag_value=0;
            end
    11824 : begin
              real_value= 0;
              imag_value=0;
            end
    11825 : begin
              real_value= 0;
              imag_value=0;
            end
    11826 : begin
              real_value= 0;
              imag_value=0;
            end
    11827 : begin
              real_value= 0;
              imag_value=0;
            end
    11828 : begin
              real_value= 0;
              imag_value=0;
            end
    11829 : begin
              real_value= 0;
              imag_value=0;
            end
    11830 : begin
              real_value= 0;
              imag_value=0;
            end
    11831 : begin
              real_value= 0;
              imag_value=0;
            end
    11832 : begin
              real_value= 0;
              imag_value=0;
            end
    11833 : begin
              real_value= 0;
              imag_value=0;
            end
    11834 : begin
              real_value= 0;
              imag_value=0;
            end
    11835 : begin
              real_value= 0;
              imag_value=0;
            end
    11836 : begin
              real_value= 0;
              imag_value=0;
            end
    11837 : begin
              real_value= 0;
              imag_value=0;
            end
    11838 : begin
              real_value= 0;
              imag_value=0;
            end
    11839 : begin
              real_value= 0;
              imag_value=0;
            end
    11840 : begin
              real_value= 0;
              imag_value=0;
            end
    11841 : begin
              real_value= 0;
              imag_value=0;
            end
    11842 : begin
              real_value= 0;
              imag_value=0;
            end
    11843 : begin
              real_value= 0;
              imag_value=0;
            end
    11844 : begin
              real_value= 0;
              imag_value=0;
            end
    11845 : begin
              real_value= 0;
              imag_value=0;
            end
    11846 : begin
              real_value= 0;
              imag_value=0;
            end
    11847 : begin
              real_value= 0;
              imag_value=0;
            end
    11848 : begin
              real_value= 0;
              imag_value=0;
            end
    11849 : begin
              real_value= 0;
              imag_value=0;
            end
    11850 : begin
              real_value= 0;
              imag_value=0;
            end
    11851 : begin
              real_value= 0;
              imag_value=0;
            end
    11852 : begin
              real_value= 0;
              imag_value=0;
            end
    11853 : begin
              real_value= 0;
              imag_value=0;
            end
    11854 : begin
              real_value= 0;
              imag_value=0;
            end
    11855 : begin
              real_value= 0;
              imag_value=0;
            end
    11856 : begin
              real_value= 0;
              imag_value=0;
            end
    11857 : begin
              real_value= 0;
              imag_value=0;
            end
    11858 : begin
              real_value= 0;
              imag_value=0;
            end
    11859 : begin
              real_value= 0;
              imag_value=0;
            end
    11860 : begin
              real_value= 0;
              imag_value=0;
            end
    11861 : begin
              real_value= 0;
              imag_value=0;
            end
    11862 : begin
              real_value= 0;
              imag_value=0;
            end
    11863 : begin
              real_value= 0;
              imag_value=0;
            end
    11864 : begin
              real_value= 0;
              imag_value=0;
            end
    11865 : begin
              real_value= 0;
              imag_value=0;
            end
    11866 : begin
              real_value= 0;
              imag_value=0;
            end
    11867 : begin
              real_value= 0;
              imag_value=0;
            end
    11868 : begin
              real_value= 0;
              imag_value=0;
            end
    11869 : begin
              real_value= 0;
              imag_value=0;
            end
    11870 : begin
              real_value= 0;
              imag_value=0;
            end
    11871 : begin
              real_value= 0;
              imag_value=0;
            end
    11872 : begin
              real_value= 0;
              imag_value=0;
            end
    11873 : begin
              real_value= 0;
              imag_value=0;
            end
    11874 : begin
              real_value= 0;
              imag_value=0;
            end
    11875 : begin
              real_value= 0;
              imag_value=0;
            end
    11876 : begin
              real_value= 0;
              imag_value=0;
            end
    11877 : begin
              real_value= 0;
              imag_value=0;
            end
    11878 : begin
              real_value= 0;
              imag_value=0;
            end
    11879 : begin
              real_value= 0;
              imag_value=0;
            end
    11880 : begin
              real_value= 0;
              imag_value=0;
            end
    11881 : begin
              real_value= 0;
              imag_value=0;
            end
    11882 : begin
              real_value= 0;
              imag_value=0;
            end
    11883 : begin
              real_value= 0;
              imag_value=0;
            end
    11884 : begin
              real_value= 0;
              imag_value=0;
            end
    11885 : begin
              real_value= 0;
              imag_value=0;
            end
    11886 : begin
              real_value= 0;
              imag_value=0;
            end
    11887 : begin
              real_value= 0;
              imag_value=0;
            end
    11888 : begin
              real_value= 0;
              imag_value=0;
            end
    11889 : begin
              real_value= 0;
              imag_value=0;
            end
    11890 : begin
              real_value= 0;
              imag_value=0;
            end
    11891 : begin
              real_value= 0;
              imag_value=0;
            end
    11892 : begin
              real_value= 0;
              imag_value=0;
            end
    11893 : begin
              real_value= 0;
              imag_value=0;
            end
    11894 : begin
              real_value= 0;
              imag_value=0;
            end
    11895 : begin
              real_value= 0;
              imag_value=0;
            end
    11896 : begin
              real_value= 0;
              imag_value=0;
            end
    11897 : begin
              real_value= 0;
              imag_value=0;
            end
    11898 : begin
              real_value= 0;
              imag_value=0;
            end
    11899 : begin
              real_value= 0;
              imag_value=0;
            end
    11900 : begin
              real_value= 0;
              imag_value=0;
            end
    11901 : begin
              real_value= 0;
              imag_value=0;
            end
    11902 : begin
              real_value= 0;
              imag_value=0;
            end
    11903 : begin
              real_value= 0;
              imag_value=0;
            end
    11904 : begin
              real_value= 0;
              imag_value=0;
            end
    11905 : begin
              real_value= 0;
              imag_value=0;
            end
    11906 : begin
              real_value= 0;
              imag_value=0;
            end
    11907 : begin
              real_value= 0;
              imag_value=0;
            end
    11908 : begin
              real_value= 0;
              imag_value=0;
            end
    11909 : begin
              real_value= 0;
              imag_value=0;
            end
    11910 : begin
              real_value= 0;
              imag_value=0;
            end
    11911 : begin
              real_value= 0;
              imag_value=0;
            end
    11912 : begin
              real_value= 0;
              imag_value=0;
            end
    11913 : begin
              real_value= 0;
              imag_value=0;
            end
    11914 : begin
              real_value= 0;
              imag_value=0;
            end
    11915 : begin
              real_value= 0;
              imag_value=0;
            end
    11916 : begin
              real_value= 0;
              imag_value=0;
            end
    11917 : begin
              real_value= 0;
              imag_value=0;
            end
    11918 : begin
              real_value= 0;
              imag_value=0;
            end
    11919 : begin
              real_value= 0;
              imag_value=0;
            end
    11920 : begin
              real_value= 0;
              imag_value=0;
            end
    11921 : begin
              real_value= 0;
              imag_value=0;
            end
    11922 : begin
              real_value= 0;
              imag_value=0;
            end
    11923 : begin
              real_value= 0;
              imag_value=0;
            end
    11924 : begin
              real_value= 0;
              imag_value=0;
            end
    11925 : begin
              real_value= 0;
              imag_value=0;
            end
    11926 : begin
              real_value= 0;
              imag_value=0;
            end
    11927 : begin
              real_value= 0;
              imag_value=0;
            end
    11928 : begin
              real_value= 0;
              imag_value=0;
            end
    11929 : begin
              real_value= 0;
              imag_value=0;
            end
    11930 : begin
              real_value= 0;
              imag_value=0;
            end
    11931 : begin
              real_value= 0;
              imag_value=0;
            end
    11932 : begin
              real_value= 0;
              imag_value=0;
            end
    11933 : begin
              real_value= 0;
              imag_value=0;
            end
    11934 : begin
              real_value= 0;
              imag_value=0;
            end
    11935 : begin
              real_value= 0;
              imag_value=0;
            end
    11936 : begin
              real_value= 0;
              imag_value=0;
            end
    11937 : begin
              real_value= 0;
              imag_value=0;
            end
    11938 : begin
              real_value= 0;
              imag_value=0;
            end
    11939 : begin
              real_value= 0;
              imag_value=0;
            end
    11940 : begin
              real_value= 0;
              imag_value=0;
            end
    11941 : begin
              real_value= 0;
              imag_value=0;
            end
    11942 : begin
              real_value= 0;
              imag_value=0;
            end
    11943 : begin
              real_value= 0;
              imag_value=0;
            end
    11944 : begin
              real_value= 0;
              imag_value=0;
            end
    11945 : begin
              real_value= 0;
              imag_value=0;
            end
    11946 : begin
              real_value= 0;
              imag_value=0;
            end
    11947 : begin
              real_value= 0;
              imag_value=0;
            end
    11948 : begin
              real_value= 0;
              imag_value=0;
            end
    11949 : begin
              real_value= 0;
              imag_value=0;
            end
    11950 : begin
              real_value= 0;
              imag_value=0;
            end
    11951 : begin
              real_value= 0;
              imag_value=0;
            end
    11952 : begin
              real_value= 0;
              imag_value=0;
            end
    11953 : begin
              real_value= 0;
              imag_value=0;
            end
    11954 : begin
              real_value= 0;
              imag_value=0;
            end
    11955 : begin
              real_value= 0;
              imag_value=0;
            end
    11956 : begin
              real_value= 0;
              imag_value=0;
            end
    11957 : begin
              real_value= 0;
              imag_value=0;
            end
    11958 : begin
              real_value= 0;
              imag_value=0;
            end
    11959 : begin
              real_value= 0;
              imag_value=0;
            end
    11960 : begin
              real_value= 0;
              imag_value=0;
            end
    11961 : begin
              real_value= 0;
              imag_value=0;
            end
    11962 : begin
              real_value= 0;
              imag_value=0;
            end
    11963 : begin
              real_value= 0;
              imag_value=0;
            end
    11964 : begin
              real_value= 0;
              imag_value=0;
            end
    11965 : begin
              real_value= 0;
              imag_value=0;
            end
    11966 : begin
              real_value= 0;
              imag_value=0;
            end
    11967 : begin
              real_value= 0;
              imag_value=0;
            end
    11968 : begin
              real_value= 0;
              imag_value=0;
            end
    11969 : begin
              real_value= 0;
              imag_value=0;
            end
    11970 : begin
              real_value= 0;
              imag_value=0;
            end
    11971 : begin
              real_value= 0;
              imag_value=0;
            end
    11972 : begin
              real_value= 0;
              imag_value=0;
            end
    11973 : begin
              real_value= 0;
              imag_value=0;
            end
    11974 : begin
              real_value= 0;
              imag_value=0;
            end
    11975 : begin
              real_value= 0;
              imag_value=0;
            end
    11976 : begin
              real_value= 0;
              imag_value=0;
            end
    11977 : begin
              real_value= 0;
              imag_value=0;
            end
    11978 : begin
              real_value= 0;
              imag_value=0;
            end
    11979 : begin
              real_value= 0;
              imag_value=0;
            end
    11980 : begin
              real_value= 0;
              imag_value=0;
            end
    11981 : begin
              real_value= 0;
              imag_value=0;
            end
    11982 : begin
              real_value= 0;
              imag_value=0;
            end
    11983 : begin
              real_value= 0;
              imag_value=0;
            end
    11984 : begin
              real_value= 0;
              imag_value=0;
            end
    11985 : begin
              real_value= 0;
              imag_value=0;
            end
    11986 : begin
              real_value= 0;
              imag_value=0;
            end
    11987 : begin
              real_value= 0;
              imag_value=0;
            end
    11988 : begin
              real_value= 0;
              imag_value=0;
            end
    11989 : begin
              real_value= 0;
              imag_value=0;
            end
    11990 : begin
              real_value= 0;
              imag_value=0;
            end
    11991 : begin
              real_value= 0;
              imag_value=0;
            end
    11992 : begin
              real_value= 0;
              imag_value=0;
            end
    11993 : begin
              real_value= 0;
              imag_value=0;
            end
    11994 : begin
              real_value= 0;
              imag_value=0;
            end
    11995 : begin
              real_value= 0;
              imag_value=0;
            end
    11996 : begin
              real_value= 0;
              imag_value=0;
            end
    11997 : begin
              real_value= 0;
              imag_value=0;
            end
    11998 : begin
              real_value= 0;
              imag_value=0;
            end
    11999 : begin
              real_value= 0;
              imag_value=0;
            end
    12000 : begin
              real_value= 0;
              imag_value=0;
            end
    12001 : begin
              real_value= 0;
              imag_value=0;
            end
    12002 : begin
              real_value= 0;
              imag_value=0;
            end
    12003 : begin
              real_value= 0;
              imag_value=0;
            end
    12004 : begin
              real_value= 0;
              imag_value=0;
            end
    12005 : begin
              real_value= 0;
              imag_value=0;
            end
    12006 : begin
              real_value= 0;
              imag_value=0;
            end
    12007 : begin
              real_value= 0;
              imag_value=0;
            end
    12008 : begin
              real_value= 0;
              imag_value=0;
            end
    12009 : begin
              real_value= 0;
              imag_value=0;
            end
    12010 : begin
              real_value= 0;
              imag_value=0;
            end
    12011 : begin
              real_value= 0;
              imag_value=0;
            end
    12012 : begin
              real_value= 0;
              imag_value=0;
            end
    12013 : begin
              real_value= 0;
              imag_value=0;
            end
    12014 : begin
              real_value= 0;
              imag_value=0;
            end
    12015 : begin
              real_value= 0;
              imag_value=0;
            end
    12016 : begin
              real_value= 0;
              imag_value=0;
            end
    12017 : begin
              real_value= 0;
              imag_value=0;
            end
    12018 : begin
              real_value= 0;
              imag_value=0;
            end
    12019 : begin
              real_value= 0;
              imag_value=0;
            end
    12020 : begin
              real_value= 0;
              imag_value=0;
            end
    12021 : begin
              real_value= 0;
              imag_value=0;
            end
    12022 : begin
              real_value= 0;
              imag_value=0;
            end
    12023 : begin
              real_value= 0;
              imag_value=0;
            end
    12024 : begin
              real_value= 0;
              imag_value=0;
            end
    12025 : begin
              real_value= 0;
              imag_value=0;
            end
    12026 : begin
              real_value= 0;
              imag_value=0;
            end
    12027 : begin
              real_value= 0;
              imag_value=0;
            end
    12028 : begin
              real_value= 0;
              imag_value=0;
            end
    12029 : begin
              real_value= 0;
              imag_value=0;
            end
    12030 : begin
              real_value= 0;
              imag_value=0;
            end
    12031 : begin
              real_value= 0;
              imag_value=0;
            end
    12032 : begin
              real_value= 0;
              imag_value=0;
            end
    12033 : begin
              real_value= 0;
              imag_value=0;
            end
    12034 : begin
              real_value= 0;
              imag_value=0;
            end
    12035 : begin
              real_value= 0;
              imag_value=0;
            end
    12036 : begin
              real_value= 0;
              imag_value=0;
            end
    12037 : begin
              real_value= 0;
              imag_value=0;
            end
    12038 : begin
              real_value= 0;
              imag_value=0;
            end
    12039 : begin
              real_value= 0;
              imag_value=0;
            end
    12040 : begin
              real_value= 0;
              imag_value=0;
            end
    12041 : begin
              real_value= 0;
              imag_value=0;
            end
    12042 : begin
              real_value= 0;
              imag_value=0;
            end
    12043 : begin
              real_value= 0;
              imag_value=0;
            end
    12044 : begin
              real_value= 0;
              imag_value=0;
            end
    12045 : begin
              real_value= 0;
              imag_value=0;
            end
    12046 : begin
              real_value= 0;
              imag_value=0;
            end
    12047 : begin
              real_value= 0;
              imag_value=0;
            end
    12048 : begin
              real_value= 0;
              imag_value=0;
            end
    12049 : begin
              real_value= 0;
              imag_value=0;
            end
    12050 : begin
              real_value= 0;
              imag_value=0;
            end
    12051 : begin
              real_value= 0;
              imag_value=0;
            end
    12052 : begin
              real_value= 0;
              imag_value=0;
            end
    12053 : begin
              real_value= 0;
              imag_value=0;
            end
    12054 : begin
              real_value= 0;
              imag_value=0;
            end
    12055 : begin
              real_value= 0;
              imag_value=0;
            end
    12056 : begin
              real_value= 0;
              imag_value=0;
            end
    12057 : begin
              real_value= 0;
              imag_value=0;
            end
    12058 : begin
              real_value= 0;
              imag_value=0;
            end
    12059 : begin
              real_value= 0;
              imag_value=0;
            end
    12060 : begin
              real_value= 0;
              imag_value=0;
            end
    12061 : begin
              real_value= 0;
              imag_value=0;
            end
    12062 : begin
              real_value= 0;
              imag_value=0;
            end
    12063 : begin
              real_value= 0;
              imag_value=0;
            end
    12064 : begin
              real_value= 0;
              imag_value=0;
            end
    12065 : begin
              real_value= 0;
              imag_value=0;
            end
    12066 : begin
              real_value= 0;
              imag_value=0;
            end
    12067 : begin
              real_value= 0;
              imag_value=0;
            end
    12068 : begin
              real_value= 0;
              imag_value=0;
            end
    12069 : begin
              real_value= 0;
              imag_value=0;
            end
    12070 : begin
              real_value= 0;
              imag_value=0;
            end
    12071 : begin
              real_value= 0;
              imag_value=0;
            end
    12072 : begin
              real_value= 0;
              imag_value=0;
            end
    12073 : begin
              real_value= 0;
              imag_value=0;
            end
    12074 : begin
              real_value= 0;
              imag_value=0;
            end
    12075 : begin
              real_value= 0;
              imag_value=0;
            end
    12076 : begin
              real_value= 0;
              imag_value=0;
            end
    12077 : begin
              real_value= 0;
              imag_value=0;
            end
    12078 : begin
              real_value= 0;
              imag_value=0;
            end
    12079 : begin
              real_value= 0;
              imag_value=0;
            end
    12080 : begin
              real_value= 0;
              imag_value=0;
            end
    12081 : begin
              real_value= 0;
              imag_value=0;
            end
    12082 : begin
              real_value= 0;
              imag_value=0;
            end
    12083 : begin
              real_value= 0;
              imag_value=0;
            end
    12084 : begin
              real_value= 0;
              imag_value=0;
            end
    12085 : begin
              real_value= 0;
              imag_value=0;
            end
    12086 : begin
              real_value= 0;
              imag_value=0;
            end
    12087 : begin
              real_value= 0;
              imag_value=0;
            end
    12088 : begin
              real_value= 0;
              imag_value=0;
            end
    12089 : begin
              real_value= 0;
              imag_value=0;
            end
    12090 : begin
              real_value= 0;
              imag_value=0;
            end
    12091 : begin
              real_value= 0;
              imag_value=0;
            end
    12092 : begin
              real_value= 0;
              imag_value=0;
            end
    12093 : begin
              real_value= 0;
              imag_value=0;
            end
    12094 : begin
              real_value= 0;
              imag_value=0;
            end
    12095 : begin
              real_value= 0;
              imag_value=0;
            end
    12096 : begin
              real_value= 0;
              imag_value=0;
            end
    12097 : begin
              real_value= 0;
              imag_value=0;
            end
    12098 : begin
              real_value= 0;
              imag_value=0;
            end
    12099 : begin
              real_value= 0;
              imag_value=0;
            end
    12100 : begin
              real_value= 0;
              imag_value=0;
            end
    12101 : begin
              real_value= 0;
              imag_value=0;
            end
    12102 : begin
              real_value= 0;
              imag_value=0;
            end
    12103 : begin
              real_value= 0;
              imag_value=0;
            end
    12104 : begin
              real_value= 0;
              imag_value=0;
            end
    12105 : begin
              real_value= 0;
              imag_value=0;
            end
    12106 : begin
              real_value= 0;
              imag_value=0;
            end
    12107 : begin
              real_value= 0;
              imag_value=0;
            end
    12108 : begin
              real_value= 0;
              imag_value=0;
            end
    12109 : begin
              real_value= 0;
              imag_value=0;
            end
    12110 : begin
              real_value= 0;
              imag_value=0;
            end
    12111 : begin
              real_value= 0;
              imag_value=0;
            end
    12112 : begin
              real_value= 0;
              imag_value=0;
            end
    12113 : begin
              real_value= 0;
              imag_value=0;
            end
    12114 : begin
              real_value= 0;
              imag_value=0;
            end
    12115 : begin
              real_value= 0;
              imag_value=0;
            end
    12116 : begin
              real_value= 0;
              imag_value=0;
            end
    12117 : begin
              real_value= 0;
              imag_value=0;
            end
    12118 : begin
              real_value= 0;
              imag_value=0;
            end
    12119 : begin
              real_value= 0;
              imag_value=0;
            end
    12120 : begin
              real_value= 0;
              imag_value=0;
            end
    12121 : begin
              real_value= 0;
              imag_value=0;
            end
    12122 : begin
              real_value= 0;
              imag_value=0;
            end
    12123 : begin
              real_value= 0;
              imag_value=0;
            end
    12124 : begin
              real_value= 0;
              imag_value=0;
            end
    12125 : begin
              real_value= 0;
              imag_value=0;
            end
    12126 : begin
              real_value= 0;
              imag_value=0;
            end
    12127 : begin
              real_value= 0;
              imag_value=0;
            end
    12128 : begin
              real_value= 0;
              imag_value=0;
            end
    12129 : begin
              real_value= 0;
              imag_value=0;
            end
    12130 : begin
              real_value= 0;
              imag_value=0;
            end
    12131 : begin
              real_value= 0;
              imag_value=0;
            end
    12132 : begin
              real_value= 0;
              imag_value=0;
            end
    12133 : begin
              real_value= 0;
              imag_value=0;
            end
    12134 : begin
              real_value= 0;
              imag_value=0;
            end
    12135 : begin
              real_value= 0;
              imag_value=0;
            end
    12136 : begin
              real_value= 0;
              imag_value=0;
            end
    12137 : begin
              real_value= 0;
              imag_value=0;
            end
    12138 : begin
              real_value= 0;
              imag_value=0;
            end
    12139 : begin
              real_value= 0;
              imag_value=0;
            end
    12140 : begin
              real_value= 0;
              imag_value=0;
            end
    12141 : begin
              real_value= 0;
              imag_value=0;
            end
    12142 : begin
              real_value= 0;
              imag_value=0;
            end
    12143 : begin
              real_value= 0;
              imag_value=0;
            end
    12144 : begin
              real_value= 0;
              imag_value=0;
            end
    12145 : begin
              real_value= 0;
              imag_value=0;
            end
    12146 : begin
              real_value= 0;
              imag_value=0;
            end
    12147 : begin
              real_value= 0;
              imag_value=0;
            end
    12148 : begin
              real_value= 0;
              imag_value=0;
            end
    12149 : begin
              real_value= 0;
              imag_value=0;
            end
    12150 : begin
              real_value= 0;
              imag_value=0;
            end
    12151 : begin
              real_value= 0;
              imag_value=0;
            end
    12152 : begin
              real_value= 0;
              imag_value=0;
            end
    12153 : begin
              real_value= 0;
              imag_value=0;
            end
    12154 : begin
              real_value= 0;
              imag_value=0;
            end
    12155 : begin
              real_value= 0;
              imag_value=0;
            end
    12156 : begin
              real_value= 0;
              imag_value=0;
            end
    12157 : begin
              real_value= 0;
              imag_value=0;
            end
    12158 : begin
              real_value= 0;
              imag_value=0;
            end
    12159 : begin
              real_value= 0;
              imag_value=0;
            end
    12160 : begin
              real_value= 0;
              imag_value=0;
            end
    12161 : begin
              real_value= 0;
              imag_value=0;
            end
    12162 : begin
              real_value= 0;
              imag_value=0;
            end
    12163 : begin
              real_value= 0;
              imag_value=0;
            end
    12164 : begin
              real_value= 0;
              imag_value=0;
            end
    12165 : begin
              real_value= 0;
              imag_value=0;
            end
    12166 : begin
              real_value= 0;
              imag_value=0;
            end
    12167 : begin
              real_value= 0;
              imag_value=0;
            end
    12168 : begin
              real_value= 0;
              imag_value=0;
            end
    12169 : begin
              real_value= 0;
              imag_value=0;
            end
    12170 : begin
              real_value= 0;
              imag_value=0;
            end
    12171 : begin
              real_value= 0;
              imag_value=0;
            end
    12172 : begin
              real_value= 0;
              imag_value=0;
            end
    12173 : begin
              real_value= 0;
              imag_value=0;
            end
    12174 : begin
              real_value= 0;
              imag_value=0;
            end
    12175 : begin
              real_value= 0;
              imag_value=0;
            end
    12176 : begin
              real_value= 0;
              imag_value=0;
            end
    12177 : begin
              real_value= 0;
              imag_value=0;
            end
    12178 : begin
              real_value= 0;
              imag_value=0;
            end
    12179 : begin
              real_value= 0;
              imag_value=0;
            end
    12180 : begin
              real_value= 0;
              imag_value=0;
            end
    12181 : begin
              real_value= 0;
              imag_value=0;
            end
    12182 : begin
              real_value= 0;
              imag_value=0;
            end
    12183 : begin
              real_value= 0;
              imag_value=0;
            end
    12184 : begin
              real_value= 0;
              imag_value=0;
            end
    12185 : begin
              real_value= 0;
              imag_value=0;
            end
    12186 : begin
              real_value= 0;
              imag_value=0;
            end
    12187 : begin
              real_value= 0;
              imag_value=0;
            end
    12188 : begin
              real_value= 0;
              imag_value=0;
            end
    12189 : begin
              real_value= 0;
              imag_value=0;
            end
    12190 : begin
              real_value= 0;
              imag_value=0;
            end
    12191 : begin
              real_value= 0;
              imag_value=0;
            end
    12192 : begin
              real_value= 0;
              imag_value=0;
            end
    12193 : begin
              real_value= 0;
              imag_value=0;
            end
    12194 : begin
              real_value= 0;
              imag_value=0;
            end
    12195 : begin
              real_value= 0;
              imag_value=0;
            end
    12196 : begin
              real_value= 0;
              imag_value=0;
            end
    12197 : begin
              real_value= 0;
              imag_value=0;
            end
    12198 : begin
              real_value= 0;
              imag_value=0;
            end
    12199 : begin
              real_value= 0;
              imag_value=0;
            end
    12200 : begin
              real_value= 0;
              imag_value=0;
            end
    12201 : begin
              real_value= 0;
              imag_value=0;
            end
    12202 : begin
              real_value= 0;
              imag_value=0;
            end
    12203 : begin
              real_value= 0;
              imag_value=0;
            end
    12204 : begin
              real_value= 0;
              imag_value=0;
            end
    12205 : begin
              real_value= 0;
              imag_value=0;
            end
    12206 : begin
              real_value= 0;
              imag_value=0;
            end
    12207 : begin
              real_value= 0;
              imag_value=0;
            end
    12208 : begin
              real_value= 0;
              imag_value=0;
            end
    12209 : begin
              real_value= 0;
              imag_value=0;
            end
    12210 : begin
              real_value= 0;
              imag_value=0;
            end
    12211 : begin
              real_value= 0;
              imag_value=0;
            end
    12212 : begin
              real_value= 0;
              imag_value=0;
            end
    12213 : begin
              real_value= 0;
              imag_value=0;
            end
    12214 : begin
              real_value= 0;
              imag_value=0;
            end
    12215 : begin
              real_value= 0;
              imag_value=0;
            end
    12216 : begin
              real_value= 0;
              imag_value=0;
            end
    12217 : begin
              real_value= 0;
              imag_value=0;
            end
    12218 : begin
              real_value= 0;
              imag_value=0;
            end
    12219 : begin
              real_value= 0;
              imag_value=0;
            end
    12220 : begin
              real_value= 0;
              imag_value=0;
            end
    12221 : begin
              real_value= 0;
              imag_value=0;
            end
    12222 : begin
              real_value= 0;
              imag_value=0;
            end
    12223 : begin
              real_value= 0;
              imag_value=0;
            end
    12224 : begin
              real_value= 0;
              imag_value=0;
            end
    12225 : begin
              real_value= 0;
              imag_value=0;
            end
    12226 : begin
              real_value= 0;
              imag_value=0;
            end
    12227 : begin
              real_value= 0;
              imag_value=0;
            end
    12228 : begin
              real_value= 0;
              imag_value=0;
            end
    12229 : begin
              real_value= 0;
              imag_value=0;
            end
    12230 : begin
              real_value= 0;
              imag_value=0;
            end
    12231 : begin
              real_value= 0;
              imag_value=0;
            end
    12232 : begin
              real_value= 0;
              imag_value=0;
            end
    12233 : begin
              real_value= 0;
              imag_value=0;
            end
    12234 : begin
              real_value= 0;
              imag_value=0;
            end
    12235 : begin
              real_value= 0;
              imag_value=0;
            end
    12236 : begin
              real_value= 0;
              imag_value=0;
            end
    12237 : begin
              real_value= 0;
              imag_value=0;
            end
    12238 : begin
              real_value= 0;
              imag_value=0;
            end
    12239 : begin
              real_value= 0;
              imag_value=0;
            end
    12240 : begin
              real_value= 0;
              imag_value=0;
            end
    12241 : begin
              real_value= 0;
              imag_value=0;
            end
    12242 : begin
              real_value= 0;
              imag_value=0;
            end
    12243 : begin
              real_value= 0;
              imag_value=0;
            end
    12244 : begin
              real_value= 0;
              imag_value=0;
            end
    12245 : begin
              real_value= 0;
              imag_value=0;
            end
    12246 : begin
              real_value= 0;
              imag_value=0;
            end
    12247 : begin
              real_value= 0;
              imag_value=0;
            end
    12248 : begin
              real_value= 0;
              imag_value=0;
            end
    12249 : begin
              real_value= 0;
              imag_value=0;
            end
    12250 : begin
              real_value= 0;
              imag_value=0;
            end
    12251 : begin
              real_value= 0;
              imag_value=0;
            end
    12252 : begin
              real_value= 0;
              imag_value=0;
            end
    12253 : begin
              real_value= 0;
              imag_value=0;
            end
    12254 : begin
              real_value= 0;
              imag_value=0;
            end
    12255 : begin
              real_value= 0;
              imag_value=0;
            end
    12256 : begin
              real_value= 0;
              imag_value=0;
            end
    12257 : begin
              real_value= 0;
              imag_value=0;
            end
    12258 : begin
              real_value= 0;
              imag_value=0;
            end
    12259 : begin
              real_value= 0;
              imag_value=0;
            end
    12260 : begin
              real_value= 0;
              imag_value=0;
            end
    12261 : begin
              real_value= 0;
              imag_value=0;
            end
    12262 : begin
              real_value= 0;
              imag_value=0;
            end
    12263 : begin
              real_value= 0;
              imag_value=0;
            end
    12264 : begin
              real_value= 0;
              imag_value=0;
            end
    12265 : begin
              real_value= 0;
              imag_value=0;
            end
    12266 : begin
              real_value= 0;
              imag_value=0;
            end
    12267 : begin
              real_value= 0;
              imag_value=0;
            end
    12268 : begin
              real_value= 0;
              imag_value=0;
            end
    12269 : begin
              real_value= 0;
              imag_value=0;
            end
    12270 : begin
              real_value= 0;
              imag_value=0;
            end
    12271 : begin
              real_value= 0;
              imag_value=0;
            end
    12272 : begin
              real_value= 0;
              imag_value=0;
            end
    12273 : begin
              real_value= 0;
              imag_value=0;
            end
    12274 : begin
              real_value= 0;
              imag_value=0;
            end
    12275 : begin
              real_value= 0;
              imag_value=0;
            end
    12276 : begin
              real_value= 0;
              imag_value=0;
            end
    12277 : begin
              real_value= 0;
              imag_value=0;
            end
    12278 : begin
              real_value= 0;
              imag_value=0;
            end
    12279 : begin
              real_value= 0;
              imag_value=0;
            end
    12280 : begin
              real_value= 0;
              imag_value=0;
            end
    12281 : begin
              real_value= 0;
              imag_value=0;
            end
    12282 : begin
              real_value= 0;
              imag_value=0;
            end
    12283 : begin
              real_value= 0;
              imag_value=0;
            end
    12284 : begin
              real_value= 0;
              imag_value=0;
            end
    12285 : begin
              real_value= 0;
              imag_value=0;
            end
    12286 : begin
              real_value= 0;
              imag_value=0;
            end
    12287 : begin
              real_value= 0;
              imag_value=0;
            end
    12288 : begin
              real_value= 0;
              imag_value=0;
            end
    12289 : begin
              real_value= 0;
              imag_value=0;
            end
    12290 : begin
              real_value= 0;
              imag_value=0;
            end
    12291 : begin
              real_value= 0;
              imag_value=0;
            end
    12292 : begin
              real_value= 0;
              imag_value=0;
            end
    12293 : begin
              real_value= 0;
              imag_value=0;
            end
    12294 : begin
              real_value= 0;
              imag_value=0;
            end
    12295 : begin
              real_value= 0;
              imag_value=0;
            end
    12296 : begin
              real_value= 0;
              imag_value=0;
            end
    12297 : begin
              real_value= 0;
              imag_value=0;
            end
    12298 : begin
              real_value= 0;
              imag_value=0;
            end
    12299 : begin
              real_value= 0;
              imag_value=0;
            end
    12300 : begin
              real_value= 0;
              imag_value=0;
            end
    12301 : begin
              real_value= 0;
              imag_value=0;
            end
    12302 : begin
              real_value= 0;
              imag_value=0;
            end
    12303 : begin
              real_value= 0;
              imag_value=0;
            end
    12304 : begin
              real_value= 0;
              imag_value=0;
            end
    12305 : begin
              real_value= 0;
              imag_value=0;
            end
    12306 : begin
              real_value= 0;
              imag_value=0;
            end
    12307 : begin
              real_value= 0;
              imag_value=0;
            end
    12308 : begin
              real_value= 0;
              imag_value=0;
            end
    12309 : begin
              real_value= 0;
              imag_value=0;
            end
    12310 : begin
              real_value= 0;
              imag_value=0;
            end
    12311 : begin
              real_value= 0;
              imag_value=0;
            end
    12312 : begin
              real_value= 0;
              imag_value=0;
            end
    12313 : begin
              real_value= 0;
              imag_value=0;
            end
    12314 : begin
              real_value= 0;
              imag_value=0;
            end
    12315 : begin
              real_value= 0;
              imag_value=0;
            end
    12316 : begin
              real_value= 0;
              imag_value=0;
            end
    12317 : begin
              real_value= 0;
              imag_value=0;
            end
    12318 : begin
              real_value= 0;
              imag_value=0;
            end
    12319 : begin
              real_value= 0;
              imag_value=0;
            end
    12320 : begin
              real_value= 0;
              imag_value=0;
            end
    12321 : begin
              real_value= 0;
              imag_value=0;
            end
    12322 : begin
              real_value= 0;
              imag_value=0;
            end
    12323 : begin
              real_value= 0;
              imag_value=0;
            end
    12324 : begin
              real_value= 0;
              imag_value=0;
            end
    12325 : begin
              real_value= 0;
              imag_value=0;
            end
    12326 : begin
              real_value= 0;
              imag_value=0;
            end
    12327 : begin
              real_value= 0;
              imag_value=0;
            end
    12328 : begin
              real_value= 0;
              imag_value=0;
            end
    12329 : begin
              real_value= 0;
              imag_value=0;
            end
    12330 : begin
              real_value= 0;
              imag_value=0;
            end
    12331 : begin
              real_value= 0;
              imag_value=0;
            end
    12332 : begin
              real_value= 0;
              imag_value=0;
            end
    12333 : begin
              real_value= 0;
              imag_value=0;
            end
    12334 : begin
              real_value= 0;
              imag_value=0;
            end
    12335 : begin
              real_value= 0;
              imag_value=0;
            end
    12336 : begin
              real_value= 0;
              imag_value=0;
            end
    12337 : begin
              real_value= 0;
              imag_value=0;
            end
    12338 : begin
              real_value= 0;
              imag_value=0;
            end
    12339 : begin
              real_value= 0;
              imag_value=0;
            end
    12340 : begin
              real_value= 0;
              imag_value=0;
            end
    12341 : begin
              real_value= 0;
              imag_value=0;
            end
    12342 : begin
              real_value= 0;
              imag_value=0;
            end
    12343 : begin
              real_value= 0;
              imag_value=0;
            end
    12344 : begin
              real_value= 0;
              imag_value=0;
            end
    12345 : begin
              real_value= 0;
              imag_value=0;
            end
    12346 : begin
              real_value= 0;
              imag_value=0;
            end
    12347 : begin
              real_value= 0;
              imag_value=0;
            end
    12348 : begin
              real_value= 0;
              imag_value=0;
            end
    12349 : begin
              real_value= 0;
              imag_value=0;
            end
    12350 : begin
              real_value= 0;
              imag_value=0;
            end
    12351 : begin
              real_value= 0;
              imag_value=0;
            end
    12352 : begin
              real_value= 0;
              imag_value=0;
            end
    12353 : begin
              real_value= 0;
              imag_value=0;
            end
    12354 : begin
              real_value= 0;
              imag_value=0;
            end
    12355 : begin
              real_value= 0;
              imag_value=0;
            end
    12356 : begin
              real_value= 0;
              imag_value=0;
            end
    12357 : begin
              real_value= 0;
              imag_value=0;
            end
    12358 : begin
              real_value= 0;
              imag_value=0;
            end
    12359 : begin
              real_value= 0;
              imag_value=0;
            end
    12360 : begin
              real_value= 0;
              imag_value=0;
            end
    12361 : begin
              real_value= 0;
              imag_value=0;
            end
    12362 : begin
              real_value= 0;
              imag_value=0;
            end
    12363 : begin
              real_value= 0;
              imag_value=0;
            end
    12364 : begin
              real_value= 0;
              imag_value=0;
            end
    12365 : begin
              real_value= 0;
              imag_value=0;
            end
    12366 : begin
              real_value= 0;
              imag_value=0;
            end
    12367 : begin
              real_value= 0;
              imag_value=0;
            end
    12368 : begin
              real_value= 0;
              imag_value=0;
            end
    12369 : begin
              real_value= 0;
              imag_value=0;
            end
    12370 : begin
              real_value= 0;
              imag_value=0;
            end
    12371 : begin
              real_value= 0;
              imag_value=0;
            end
    12372 : begin
              real_value= 0;
              imag_value=0;
            end
    12373 : begin
              real_value= 0;
              imag_value=0;
            end
    12374 : begin
              real_value= 0;
              imag_value=0;
            end
    12375 : begin
              real_value= 0;
              imag_value=0;
            end
    12376 : begin
              real_value= 0;
              imag_value=0;
            end
    12377 : begin
              real_value= 0;
              imag_value=0;
            end
    12378 : begin
              real_value= 0;
              imag_value=0;
            end
    12379 : begin
              real_value= 0;
              imag_value=0;
            end
    12380 : begin
              real_value= 0;
              imag_value=0;
            end
    12381 : begin
              real_value= 0;
              imag_value=0;
            end
    12382 : begin
              real_value= 0;
              imag_value=0;
            end
    12383 : begin
              real_value= 0;
              imag_value=0;
            end
    12384 : begin
              real_value= 0;
              imag_value=0;
            end
    12385 : begin
              real_value= 0;
              imag_value=0;
            end
    12386 : begin
              real_value= 0;
              imag_value=0;
            end
    12387 : begin
              real_value= 0;
              imag_value=0;
            end
    12388 : begin
              real_value= 0;
              imag_value=0;
            end
    12389 : begin
              real_value= 0;
              imag_value=0;
            end
    12390 : begin
              real_value= 0;
              imag_value=0;
            end
    12391 : begin
              real_value= 0;
              imag_value=0;
            end
    12392 : begin
              real_value= 0;
              imag_value=0;
            end
    12393 : begin
              real_value= 0;
              imag_value=0;
            end
    12394 : begin
              real_value= 0;
              imag_value=0;
            end
    12395 : begin
              real_value= 0;
              imag_value=0;
            end
    12396 : begin
              real_value= 0;
              imag_value=0;
            end
    12397 : begin
              real_value= 0;
              imag_value=0;
            end
    12398 : begin
              real_value= 0;
              imag_value=0;
            end
    12399 : begin
              real_value= 0;
              imag_value=0;
            end
    12400 : begin
              real_value= 0;
              imag_value=0;
            end
    12401 : begin
              real_value= 0;
              imag_value=0;
            end
    12402 : begin
              real_value= 0;
              imag_value=0;
            end
    12403 : begin
              real_value= 0;
              imag_value=0;
            end
    12404 : begin
              real_value= 0;
              imag_value=0;
            end
    12405 : begin
              real_value= 0;
              imag_value=0;
            end
    12406 : begin
              real_value= 0;
              imag_value=0;
            end
    12407 : begin
              real_value= 0;
              imag_value=0;
            end
    12408 : begin
              real_value= 0;
              imag_value=0;
            end
    12409 : begin
              real_value= 0;
              imag_value=0;
            end
    12410 : begin
              real_value= 0;
              imag_value=0;
            end
    12411 : begin
              real_value= 0;
              imag_value=0;
            end
    12412 : begin
              real_value= 0;
              imag_value=0;
            end
    12413 : begin
              real_value= 0;
              imag_value=0;
            end
    12414 : begin
              real_value= 0;
              imag_value=0;
            end
    12415 : begin
              real_value= 0;
              imag_value=0;
            end
    12416 : begin
              real_value= 0;
              imag_value=0;
            end
    12417 : begin
              real_value= 0;
              imag_value=0;
            end
    12418 : begin
              real_value= 0;
              imag_value=0;
            end
    12419 : begin
              real_value= 0;
              imag_value=0;
            end
    12420 : begin
              real_value= 0;
              imag_value=0;
            end
    12421 : begin
              real_value= 0;
              imag_value=0;
            end
    12422 : begin
              real_value= 0;
              imag_value=0;
            end
    12423 : begin
              real_value= 0;
              imag_value=0;
            end
    12424 : begin
              real_value= 0;
              imag_value=0;
            end
    12425 : begin
              real_value= 0;
              imag_value=0;
            end
    12426 : begin
              real_value= 0;
              imag_value=0;
            end
    12427 : begin
              real_value= 0;
              imag_value=0;
            end
    12428 : begin
              real_value= 0;
              imag_value=0;
            end
    12429 : begin
              real_value= 0;
              imag_value=0;
            end
    12430 : begin
              real_value= 0;
              imag_value=0;
            end
    12431 : begin
              real_value= 0;
              imag_value=0;
            end
    12432 : begin
              real_value= 0;
              imag_value=0;
            end
    12433 : begin
              real_value= 0;
              imag_value=0;
            end
    12434 : begin
              real_value= 0;
              imag_value=0;
            end
    12435 : begin
              real_value= 0;
              imag_value=0;
            end
    12436 : begin
              real_value= 0;
              imag_value=0;
            end
    12437 : begin
              real_value= 0;
              imag_value=0;
            end
    12438 : begin
              real_value= 0;
              imag_value=0;
            end
    12439 : begin
              real_value= 0;
              imag_value=0;
            end
    12440 : begin
              real_value= 0;
              imag_value=0;
            end
    12441 : begin
              real_value= 0;
              imag_value=0;
            end
    12442 : begin
              real_value= 0;
              imag_value=0;
            end
    12443 : begin
              real_value= 0;
              imag_value=0;
            end
    12444 : begin
              real_value= 0;
              imag_value=0;
            end
    12445 : begin
              real_value= 0;
              imag_value=0;
            end
    12446 : begin
              real_value= 0;
              imag_value=0;
            end
    12447 : begin
              real_value= 0;
              imag_value=0;
            end
    12448 : begin
              real_value= 0;
              imag_value=0;
            end
    12449 : begin
              real_value= 0;
              imag_value=0;
            end
    12450 : begin
              real_value= 0;
              imag_value=0;
            end
    12451 : begin
              real_value= 0;
              imag_value=0;
            end
    12452 : begin
              real_value= 0;
              imag_value=0;
            end
    12453 : begin
              real_value= 0;
              imag_value=0;
            end
    12454 : begin
              real_value= 0;
              imag_value=0;
            end
    12455 : begin
              real_value= 0;
              imag_value=0;
            end
    12456 : begin
              real_value= 0;
              imag_value=0;
            end
    12457 : begin
              real_value= 0;
              imag_value=0;
            end
    12458 : begin
              real_value= 0;
              imag_value=0;
            end
    12459 : begin
              real_value= 0;
              imag_value=0;
            end
    12460 : begin
              real_value= 0;
              imag_value=0;
            end
    12461 : begin
              real_value= 0;
              imag_value=0;
            end
    12462 : begin
              real_value= 0;
              imag_value=0;
            end
    12463 : begin
              real_value= 0;
              imag_value=0;
            end
    12464 : begin
              real_value= 0;
              imag_value=0;
            end
    12465 : begin
              real_value= 0;
              imag_value=0;
            end
    12466 : begin
              real_value= 0;
              imag_value=0;
            end
    12467 : begin
              real_value= 0;
              imag_value=0;
            end
    12468 : begin
              real_value= 0;
              imag_value=0;
            end
    12469 : begin
              real_value= 0;
              imag_value=0;
            end
    12470 : begin
              real_value= 0;
              imag_value=0;
            end
    12471 : begin
              real_value= 0;
              imag_value=0;
            end
    12472 : begin
              real_value= 0;
              imag_value=0;
            end
    12473 : begin
              real_value= 0;
              imag_value=0;
            end
    12474 : begin
              real_value= 0;
              imag_value=0;
            end
    12475 : begin
              real_value= 0;
              imag_value=0;
            end
    12476 : begin
              real_value= 0;
              imag_value=0;
            end
    12477 : begin
              real_value= 0;
              imag_value=0;
            end
    12478 : begin
              real_value= 0;
              imag_value=0;
            end
    12479 : begin
              real_value= 0;
              imag_value=0;
            end
    12480 : begin
              real_value= 0;
              imag_value=0;
            end
    12481 : begin
              real_value= 0;
              imag_value=0;
            end
    12482 : begin
              real_value= 0;
              imag_value=0;
            end
    12483 : begin
              real_value= 0;
              imag_value=0;
            end
    12484 : begin
              real_value= 0;
              imag_value=0;
            end
    12485 : begin
              real_value= 0;
              imag_value=0;
            end
    12486 : begin
              real_value= 0;
              imag_value=0;
            end
    12487 : begin
              real_value= 0;
              imag_value=0;
            end
    12488 : begin
              real_value= 0;
              imag_value=0;
            end
    12489 : begin
              real_value= 0;
              imag_value=0;
            end
    12490 : begin
              real_value= 0;
              imag_value=0;
            end
    12491 : begin
              real_value= 0;
              imag_value=0;
            end
    12492 : begin
              real_value= 0;
              imag_value=0;
            end
    12493 : begin
              real_value= 0;
              imag_value=0;
            end
    12494 : begin
              real_value= 0;
              imag_value=0;
            end
    12495 : begin
              real_value= 0;
              imag_value=0;
            end
    12496 : begin
              real_value= 0;
              imag_value=0;
            end
    12497 : begin
              real_value= 0;
              imag_value=0;
            end
    12498 : begin
              real_value= 0;
              imag_value=0;
            end
    12499 : begin
              real_value= 0;
              imag_value=0;
            end
    12500 : begin
              real_value= 0;
              imag_value=0;
            end
    12501 : begin
              real_value= 0;
              imag_value=0;
            end
    12502 : begin
              real_value= 0;
              imag_value=0;
            end
    12503 : begin
              real_value= 0;
              imag_value=0;
            end
    12504 : begin
              real_value= 0;
              imag_value=0;
            end
    12505 : begin
              real_value= 0;
              imag_value=0;
            end
    12506 : begin
              real_value= 0;
              imag_value=0;
            end
    12507 : begin
              real_value= 0;
              imag_value=0;
            end
    12508 : begin
              real_value= 0;
              imag_value=0;
            end
    12509 : begin
              real_value= 0;
              imag_value=0;
            end
    12510 : begin
              real_value= 0;
              imag_value=0;
            end
    12511 : begin
              real_value= 0;
              imag_value=0;
            end
    12512 : begin
              real_value= 0;
              imag_value=0;
            end
    12513 : begin
              real_value= 0;
              imag_value=0;
            end
    12514 : begin
              real_value= 0;
              imag_value=0;
            end
    12515 : begin
              real_value= 0;
              imag_value=0;
            end
    12516 : begin
              real_value= 0;
              imag_value=0;
            end
    12517 : begin
              real_value= 0;
              imag_value=0;
            end
    12518 : begin
              real_value= 0;
              imag_value=0;
            end
    12519 : begin
              real_value= 0;
              imag_value=0;
            end
    12520 : begin
              real_value= 0;
              imag_value=0;
            end
    12521 : begin
              real_value= 0;
              imag_value=0;
            end
    12522 : begin
              real_value= 0;
              imag_value=0;
            end
    12523 : begin
              real_value= 0;
              imag_value=0;
            end
    12524 : begin
              real_value= 0;
              imag_value=0;
            end
    12525 : begin
              real_value= 0;
              imag_value=0;
            end
    12526 : begin
              real_value= 0;
              imag_value=0;
            end
    12527 : begin
              real_value= 0;
              imag_value=0;
            end
    12528 : begin
              real_value= 0;
              imag_value=0;
            end
    12529 : begin
              real_value= 0;
              imag_value=0;
            end
    12530 : begin
              real_value= 0;
              imag_value=0;
            end
    12531 : begin
              real_value= 0;
              imag_value=0;
            end
    12532 : begin
              real_value= 0;
              imag_value=0;
            end
    12533 : begin
              real_value= 0;
              imag_value=0;
            end
    12534 : begin
              real_value= 0;
              imag_value=0;
            end
    12535 : begin
              real_value= 0;
              imag_value=0;
            end
    12536 : begin
              real_value= 0;
              imag_value=0;
            end
    12537 : begin
              real_value= 0;
              imag_value=0;
            end
    12538 : begin
              real_value= 0;
              imag_value=0;
            end
    12539 : begin
              real_value= 0;
              imag_value=0;
            end
    12540 : begin
              real_value= 0;
              imag_value=0;
            end
    12541 : begin
              real_value= 0;
              imag_value=0;
            end
    12542 : begin
              real_value= 0;
              imag_value=0;
            end
    12543 : begin
              real_value= 0;
              imag_value=0;
            end
    12544 : begin
              real_value= 0;
              imag_value=0;
            end
    12545 : begin
              real_value= 0;
              imag_value=0;
            end
    12546 : begin
              real_value= 0;
              imag_value=0;
            end
    12547 : begin
              real_value= 0;
              imag_value=0;
            end
    12548 : begin
              real_value= 0;
              imag_value=0;
            end
    12549 : begin
              real_value= 0;
              imag_value=0;
            end
    12550 : begin
              real_value= 0;
              imag_value=0;
            end
    12551 : begin
              real_value= 0;
              imag_value=0;
            end
    12552 : begin
              real_value= 0;
              imag_value=0;
            end
    12553 : begin
              real_value= 0;
              imag_value=0;
            end
    12554 : begin
              real_value= 0;
              imag_value=0;
            end
    12555 : begin
              real_value= 0;
              imag_value=0;
            end
    12556 : begin
              real_value= 0;
              imag_value=0;
            end
    12557 : begin
              real_value= 0;
              imag_value=0;
            end
    12558 : begin
              real_value= 0;
              imag_value=0;
            end
    12559 : begin
              real_value= 0;
              imag_value=0;
            end
    12560 : begin
              real_value= 0;
              imag_value=0;
            end
    12561 : begin
              real_value= 0;
              imag_value=0;
            end
    12562 : begin
              real_value= 0;
              imag_value=0;
            end
    12563 : begin
              real_value= 0;
              imag_value=0;
            end
    12564 : begin
              real_value= 0;
              imag_value=0;
            end
    12565 : begin
              real_value= 0;
              imag_value=0;
            end
    12566 : begin
              real_value= 0;
              imag_value=0;
            end
    12567 : begin
              real_value= 0;
              imag_value=0;
            end
    12568 : begin
              real_value= 0;
              imag_value=0;
            end
    12569 : begin
              real_value= 0;
              imag_value=0;
            end
    12570 : begin
              real_value= 0;
              imag_value=0;
            end
    12571 : begin
              real_value= 0;
              imag_value=0;
            end
    12572 : begin
              real_value= 0;
              imag_value=0;
            end
    12573 : begin
              real_value= 0;
              imag_value=0;
            end
    12574 : begin
              real_value= 0;
              imag_value=0;
            end
    12575 : begin
              real_value= 0;
              imag_value=0;
            end
    12576 : begin
              real_value= 0;
              imag_value=0;
            end
    12577 : begin
              real_value= 0;
              imag_value=0;
            end
    12578 : begin
              real_value= 0;
              imag_value=0;
            end
    12579 : begin
              real_value= 0;
              imag_value=0;
            end
    12580 : begin
              real_value= 0;
              imag_value=0;
            end
    12581 : begin
              real_value= 0;
              imag_value=0;
            end
    12582 : begin
              real_value= 0;
              imag_value=0;
            end
    12583 : begin
              real_value= 0;
              imag_value=0;
            end
    12584 : begin
              real_value= 0;
              imag_value=0;
            end
    12585 : begin
              real_value= 0;
              imag_value=0;
            end
    12586 : begin
              real_value= 0;
              imag_value=0;
            end
    12587 : begin
              real_value= 0;
              imag_value=0;
            end
    12588 : begin
              real_value= 0;
              imag_value=0;
            end
    12589 : begin
              real_value= 0;
              imag_value=0;
            end
    12590 : begin
              real_value= 0;
              imag_value=0;
            end
    12591 : begin
              real_value= 0;
              imag_value=0;
            end
    12592 : begin
              real_value= 0;
              imag_value=0;
            end
    12593 : begin
              real_value= 0;
              imag_value=0;
            end
    12594 : begin
              real_value= 0;
              imag_value=0;
            end
    12595 : begin
              real_value= 0;
              imag_value=0;
            end
    12596 : begin
              real_value= 0;
              imag_value=0;
            end
    12597 : begin
              real_value= 0;
              imag_value=0;
            end
    12598 : begin
              real_value= 0;
              imag_value=0;
            end
    12599 : begin
              real_value= 0;
              imag_value=0;
            end
    12600 : begin
              real_value= 0;
              imag_value=0;
            end
    12601 : begin
              real_value= 0;
              imag_value=0;
            end
    12602 : begin
              real_value= 0;
              imag_value=0;
            end
    12603 : begin
              real_value= 0;
              imag_value=0;
            end
    12604 : begin
              real_value= 0;
              imag_value=0;
            end
    12605 : begin
              real_value= 0;
              imag_value=0;
            end
    12606 : begin
              real_value= 0;
              imag_value=0;
            end
    12607 : begin
              real_value= 0;
              imag_value=0;
            end
    12608 : begin
              real_value= 0;
              imag_value=0;
            end
    12609 : begin
              real_value= 0;
              imag_value=0;
            end
    12610 : begin
              real_value= 0;
              imag_value=0;
            end
    12611 : begin
              real_value= 0;
              imag_value=0;
            end
    12612 : begin
              real_value= 0;
              imag_value=0;
            end
    12613 : begin
              real_value= 0;
              imag_value=0;
            end
    12614 : begin
              real_value= 0;
              imag_value=0;
            end
    12615 : begin
              real_value= 0;
              imag_value=0;
            end
    12616 : begin
              real_value= 0;
              imag_value=0;
            end
    12617 : begin
              real_value= 0;
              imag_value=0;
            end
    12618 : begin
              real_value= 0;
              imag_value=0;
            end
    12619 : begin
              real_value= 0;
              imag_value=0;
            end
    12620 : begin
              real_value= 0;
              imag_value=0;
            end
    12621 : begin
              real_value= 0;
              imag_value=0;
            end
    12622 : begin
              real_value= 0;
              imag_value=0;
            end
    12623 : begin
              real_value= 0;
              imag_value=0;
            end
    12624 : begin
              real_value= 0;
              imag_value=0;
            end
    12625 : begin
              real_value= 0;
              imag_value=0;
            end
    12626 : begin
              real_value= 0;
              imag_value=0;
            end
    12627 : begin
              real_value= 0;
              imag_value=0;
            end
    12628 : begin
              real_value= 0;
              imag_value=0;
            end
    12629 : begin
              real_value= 0;
              imag_value=0;
            end
    12630 : begin
              real_value= 0;
              imag_value=0;
            end
    12631 : begin
              real_value= 0;
              imag_value=0;
            end
    12632 : begin
              real_value= 0;
              imag_value=0;
            end
    12633 : begin
              real_value= 0;
              imag_value=0;
            end
    12634 : begin
              real_value= 0;
              imag_value=0;
            end
    12635 : begin
              real_value= 0;
              imag_value=0;
            end
    12636 : begin
              real_value= 0;
              imag_value=0;
            end
    12637 : begin
              real_value= 0;
              imag_value=0;
            end
    12638 : begin
              real_value= 0;
              imag_value=0;
            end
    12639 : begin
              real_value= 0;
              imag_value=0;
            end
    12640 : begin
              real_value= 0;
              imag_value=0;
            end
    12641 : begin
              real_value= 0;
              imag_value=0;
            end
    12642 : begin
              real_value= 0;
              imag_value=0;
            end
    12643 : begin
              real_value= 0;
              imag_value=0;
            end
    12644 : begin
              real_value= 0;
              imag_value=0;
            end
    12645 : begin
              real_value= 0;
              imag_value=0;
            end
    12646 : begin
              real_value= 0;
              imag_value=0;
            end
    12647 : begin
              real_value= 0;
              imag_value=0;
            end
    12648 : begin
              real_value= 0;
              imag_value=0;
            end
    12649 : begin
              real_value= 0;
              imag_value=0;
            end
    12650 : begin
              real_value= 0;
              imag_value=0;
            end
    12651 : begin
              real_value= 0;
              imag_value=0;
            end
    12652 : begin
              real_value= 0;
              imag_value=0;
            end
    12653 : begin
              real_value= 0;
              imag_value=0;
            end
    12654 : begin
              real_value= 0;
              imag_value=0;
            end
    12655 : begin
              real_value= 0;
              imag_value=0;
            end
    12656 : begin
              real_value= 0;
              imag_value=0;
            end
    12657 : begin
              real_value= 0;
              imag_value=0;
            end
    12658 : begin
              real_value= 0;
              imag_value=0;
            end
    12659 : begin
              real_value= 0;
              imag_value=0;
            end
    12660 : begin
              real_value= 0;
              imag_value=0;
            end
    12661 : begin
              real_value= 0;
              imag_value=0;
            end
    12662 : begin
              real_value= 0;
              imag_value=0;
            end
    12663 : begin
              real_value= 0;
              imag_value=0;
            end
    12664 : begin
              real_value= 0;
              imag_value=0;
            end
    12665 : begin
              real_value= 0;
              imag_value=0;
            end
    12666 : begin
              real_value= 0;
              imag_value=0;
            end
    12667 : begin
              real_value= 0;
              imag_value=0;
            end
    12668 : begin
              real_value= 0;
              imag_value=0;
            end
    12669 : begin
              real_value= 0;
              imag_value=0;
            end
    12670 : begin
              real_value= 0;
              imag_value=0;
            end
    12671 : begin
              real_value= 0;
              imag_value=0;
            end
    12672 : begin
              real_value= 0;
              imag_value=0;
            end
    12673 : begin
              real_value= 0;
              imag_value=0;
            end
    12674 : begin
              real_value= 0;
              imag_value=0;
            end
    12675 : begin
              real_value= 0;
              imag_value=0;
            end
    12676 : begin
              real_value= 0;
              imag_value=0;
            end
    12677 : begin
              real_value= 0;
              imag_value=0;
            end
    12678 : begin
              real_value= 0;
              imag_value=0;
            end
    12679 : begin
              real_value= 0;
              imag_value=0;
            end
    12680 : begin
              real_value= 0;
              imag_value=0;
            end
    12681 : begin
              real_value= 0;
              imag_value=0;
            end
    12682 : begin
              real_value= 0;
              imag_value=0;
            end
    12683 : begin
              real_value= 0;
              imag_value=0;
            end
    12684 : begin
              real_value= 0;
              imag_value=0;
            end
    12685 : begin
              real_value= 0;
              imag_value=0;
            end
    12686 : begin
              real_value= 0;
              imag_value=0;
            end
    12687 : begin
              real_value= 0;
              imag_value=0;
            end
    12688 : begin
              real_value= 0;
              imag_value=0;
            end
    12689 : begin
              real_value= 0;
              imag_value=0;
            end
    12690 : begin
              real_value= 0;
              imag_value=0;
            end
    12691 : begin
              real_value= 0;
              imag_value=0;
            end
    12692 : begin
              real_value= 0;
              imag_value=0;
            end
    12693 : begin
              real_value= 0;
              imag_value=0;
            end
    12694 : begin
              real_value= 0;
              imag_value=0;
            end
    12695 : begin
              real_value= 0;
              imag_value=0;
            end
    12696 : begin
              real_value= 0;
              imag_value=0;
            end
    12697 : begin
              real_value= 0;
              imag_value=0;
            end
    12698 : begin
              real_value= 0;
              imag_value=0;
            end
    12699 : begin
              real_value= 0;
              imag_value=0;
            end
    12700 : begin
              real_value= 0;
              imag_value=0;
            end
    12701 : begin
              real_value= 0;
              imag_value=0;
            end
    12702 : begin
              real_value= 0;
              imag_value=0;
            end
    12703 : begin
              real_value= 0;
              imag_value=0;
            end
    12704 : begin
              real_value= 0;
              imag_value=0;
            end
    12705 : begin
              real_value= 0;
              imag_value=0;
            end
    12706 : begin
              real_value= 0;
              imag_value=0;
            end
    12707 : begin
              real_value= 0;
              imag_value=0;
            end
    12708 : begin
              real_value= 0;
              imag_value=0;
            end
    12709 : begin
              real_value= 0;
              imag_value=0;
            end
    12710 : begin
              real_value= 0;
              imag_value=0;
            end
    12711 : begin
              real_value= 0;
              imag_value=0;
            end
    12712 : begin
              real_value= 0;
              imag_value=0;
            end
    12713 : begin
              real_value= 0;
              imag_value=0;
            end
    12714 : begin
              real_value= 0;
              imag_value=0;
            end
    12715 : begin
              real_value= 0;
              imag_value=0;
            end
    12716 : begin
              real_value= 0;
              imag_value=0;
            end
    12717 : begin
              real_value= 0;
              imag_value=0;
            end
    12718 : begin
              real_value= 0;
              imag_value=0;
            end
    12719 : begin
              real_value= 0;
              imag_value=0;
            end
    12720 : begin
              real_value= 0;
              imag_value=0;
            end
    12721 : begin
              real_value= 0;
              imag_value=0;
            end
    12722 : begin
              real_value= 0;
              imag_value=0;
            end
    12723 : begin
              real_value= 0;
              imag_value=0;
            end
    12724 : begin
              real_value= 0;
              imag_value=0;
            end
    12725 : begin
              real_value= 0;
              imag_value=0;
            end
    12726 : begin
              real_value= 0;
              imag_value=0;
            end
    12727 : begin
              real_value= 0;
              imag_value=0;
            end
    12728 : begin
              real_value= 0;
              imag_value=0;
            end
    12729 : begin
              real_value= 0;
              imag_value=0;
            end
    12730 : begin
              real_value= 0;
              imag_value=0;
            end
    12731 : begin
              real_value= 0;
              imag_value=0;
            end
    12732 : begin
              real_value= 0;
              imag_value=0;
            end
    12733 : begin
              real_value= 0;
              imag_value=0;
            end
    12734 : begin
              real_value= 0;
              imag_value=0;
            end
    12735 : begin
              real_value= 0;
              imag_value=0;
            end
    12736 : begin
              real_value= 0;
              imag_value=0;
            end
    12737 : begin
              real_value= 0;
              imag_value=0;
            end
    12738 : begin
              real_value= 0;
              imag_value=0;
            end
    12739 : begin
              real_value= 0;
              imag_value=0;
            end
    12740 : begin
              real_value= 0;
              imag_value=0;
            end
    12741 : begin
              real_value= 0;
              imag_value=0;
            end
    12742 : begin
              real_value= 0;
              imag_value=0;
            end
    12743 : begin
              real_value= 0;
              imag_value=0;
            end
    12744 : begin
              real_value= 0;
              imag_value=0;
            end
    12745 : begin
              real_value= 0;
              imag_value=0;
            end
    12746 : begin
              real_value= 0;
              imag_value=0;
            end
    12747 : begin
              real_value= 0;
              imag_value=0;
            end
    12748 : begin
              real_value= 0;
              imag_value=0;
            end
    12749 : begin
              real_value= 0;
              imag_value=0;
            end
    12750 : begin
              real_value= 0;
              imag_value=0;
            end
    12751 : begin
              real_value= 0;
              imag_value=0;
            end
    12752 : begin
              real_value= 0;
              imag_value=0;
            end
    12753 : begin
              real_value= 0;
              imag_value=0;
            end
    12754 : begin
              real_value= 0;
              imag_value=0;
            end
    12755 : begin
              real_value= 0;
              imag_value=0;
            end
    12756 : begin
              real_value= 0;
              imag_value=0;
            end
    12757 : begin
              real_value= 0;
              imag_value=0;
            end
    12758 : begin
              real_value= 0;
              imag_value=0;
            end
    12759 : begin
              real_value= 0;
              imag_value=0;
            end
    12760 : begin
              real_value= 0;
              imag_value=0;
            end
    12761 : begin
              real_value= 0;
              imag_value=0;
            end
    12762 : begin
              real_value= 0;
              imag_value=0;
            end
    12763 : begin
              real_value= 0;
              imag_value=0;
            end
    12764 : begin
              real_value= 0;
              imag_value=0;
            end
    12765 : begin
              real_value= 0;
              imag_value=0;
            end
    12766 : begin
              real_value= 0;
              imag_value=0;
            end
    12767 : begin
              real_value= 0;
              imag_value=0;
            end
    12768 : begin
              real_value= 0;
              imag_value=0;
            end
    12769 : begin
              real_value= 0;
              imag_value=0;
            end
    12770 : begin
              real_value= 0;
              imag_value=0;
            end
    12771 : begin
              real_value= 0;
              imag_value=0;
            end
    12772 : begin
              real_value= 0;
              imag_value=0;
            end
    12773 : begin
              real_value= 0;
              imag_value=0;
            end
    12774 : begin
              real_value= 0;
              imag_value=0;
            end
    12775 : begin
              real_value= 0;
              imag_value=0;
            end
    12776 : begin
              real_value= 0;
              imag_value=0;
            end
    12777 : begin
              real_value= 0;
              imag_value=0;
            end
    12778 : begin
              real_value= 0;
              imag_value=0;
            end
    12779 : begin
              real_value= 0;
              imag_value=0;
            end
    12780 : begin
              real_value= 0;
              imag_value=0;
            end
    12781 : begin
              real_value= 0;
              imag_value=0;
            end
    12782 : begin
              real_value= 0;
              imag_value=0;
            end
    12783 : begin
              real_value= 0;
              imag_value=0;
            end
    12784 : begin
              real_value= 0;
              imag_value=0;
            end
    12785 : begin
              real_value= 0;
              imag_value=0;
            end
    12786 : begin
              real_value= 0;
              imag_value=0;
            end
    12787 : begin
              real_value= 0;
              imag_value=0;
            end
    12788 : begin
              real_value= 0;
              imag_value=0;
            end
    12789 : begin
              real_value= 0;
              imag_value=0;
            end
    12790 : begin
              real_value= 0;
              imag_value=0;
            end
    12791 : begin
              real_value= 0;
              imag_value=0;
            end
    12792 : begin
              real_value= 0;
              imag_value=0;
            end
    12793 : begin
              real_value= 0;
              imag_value=0;
            end
    12794 : begin
              real_value= 0;
              imag_value=0;
            end
    12795 : begin
              real_value= 0;
              imag_value=0;
            end
    12796 : begin
              real_value= 0;
              imag_value=0;
            end
    12797 : begin
              real_value= 0;
              imag_value=0;
            end
    12798 : begin
              real_value= 0;
              imag_value=0;
            end
    12799 : begin
              real_value= 0;
              imag_value=0;
            end
    12800 : begin
              real_value= 0;
              imag_value=0;
            end
    12801 : begin
              real_value= 0;
              imag_value=0;
            end
    12802 : begin
              real_value= 0;
              imag_value=0;
            end
    12803 : begin
              real_value= 0;
              imag_value=0;
            end
    12804 : begin
              real_value= 0;
              imag_value=0;
            end
    12805 : begin
              real_value= 0;
              imag_value=0;
            end
    12806 : begin
              real_value= 0;
              imag_value=0;
            end
    12807 : begin
              real_value= 0;
              imag_value=0;
            end
    12808 : begin
              real_value= 0;
              imag_value=0;
            end
    12809 : begin
              real_value= 0;
              imag_value=0;
            end
    12810 : begin
              real_value= 0;
              imag_value=0;
            end
    12811 : begin
              real_value= 0;
              imag_value=0;
            end
    12812 : begin
              real_value= 0;
              imag_value=0;
            end
    12813 : begin
              real_value= 0;
              imag_value=0;
            end
    12814 : begin
              real_value= 0;
              imag_value=0;
            end
    12815 : begin
              real_value= 0;
              imag_value=0;
            end
    12816 : begin
              real_value= 0;
              imag_value=0;
            end
    12817 : begin
              real_value= 0;
              imag_value=0;
            end
    12818 : begin
              real_value= 0;
              imag_value=0;
            end
    12819 : begin
              real_value= 0;
              imag_value=0;
            end
    12820 : begin
              real_value= 0;
              imag_value=0;
            end
    12821 : begin
              real_value= 0;
              imag_value=0;
            end
    12822 : begin
              real_value= 0;
              imag_value=0;
            end
    12823 : begin
              real_value= 0;
              imag_value=0;
            end
    12824 : begin
              real_value= 0;
              imag_value=0;
            end
    12825 : begin
              real_value= 0;
              imag_value=0;
            end
    12826 : begin
              real_value= 0;
              imag_value=0;
            end
    12827 : begin
              real_value= 0;
              imag_value=0;
            end
    12828 : begin
              real_value= 0;
              imag_value=0;
            end
    12829 : begin
              real_value= 0;
              imag_value=0;
            end
    12830 : begin
              real_value= 0;
              imag_value=0;
            end
    12831 : begin
              real_value= 0;
              imag_value=0;
            end
    12832 : begin
              real_value= 0;
              imag_value=0;
            end
    12833 : begin
              real_value= 0;
              imag_value=0;
            end
    12834 : begin
              real_value= 0;
              imag_value=0;
            end
    12835 : begin
              real_value= 0;
              imag_value=0;
            end
    12836 : begin
              real_value= 0;
              imag_value=0;
            end
    12837 : begin
              real_value= 0;
              imag_value=0;
            end
    12838 : begin
              real_value= 0;
              imag_value=0;
            end
    12839 : begin
              real_value= 0;
              imag_value=0;
            end
    12840 : begin
              real_value= 0;
              imag_value=0;
            end
    12841 : begin
              real_value= 0;
              imag_value=0;
            end
    12842 : begin
              real_value= 0;
              imag_value=0;
            end
    12843 : begin
              real_value= 0;
              imag_value=0;
            end
    12844 : begin
              real_value= 0;
              imag_value=0;
            end
    12845 : begin
              real_value= 0;
              imag_value=0;
            end
    12846 : begin
              real_value= 0;
              imag_value=0;
            end
    12847 : begin
              real_value= 0;
              imag_value=0;
            end
    12848 : begin
              real_value= 0;
              imag_value=0;
            end
    12849 : begin
              real_value= 0;
              imag_value=0;
            end
    12850 : begin
              real_value= 0;
              imag_value=0;
            end
    12851 : begin
              real_value= 0;
              imag_value=0;
            end
    12852 : begin
              real_value= 0;
              imag_value=0;
            end
    12853 : begin
              real_value= 0;
              imag_value=0;
            end
    12854 : begin
              real_value= 0;
              imag_value=0;
            end
    12855 : begin
              real_value= 0;
              imag_value=0;
            end
    12856 : begin
              real_value= 0;
              imag_value=0;
            end
    12857 : begin
              real_value= 0;
              imag_value=0;
            end
    12858 : begin
              real_value= 0;
              imag_value=0;
            end
    12859 : begin
              real_value= 0;
              imag_value=0;
            end
    12860 : begin
              real_value= 0;
              imag_value=0;
            end
    12861 : begin
              real_value= 0;
              imag_value=0;
            end
    12862 : begin
              real_value= 0;
              imag_value=0;
            end
    12863 : begin
              real_value= 0;
              imag_value=0;
            end
    12864 : begin
              real_value= 0;
              imag_value=0;
            end
    12865 : begin
              real_value= 0;
              imag_value=0;
            end
    12866 : begin
              real_value= 0;
              imag_value=0;
            end
    12867 : begin
              real_value= 0;
              imag_value=0;
            end
    12868 : begin
              real_value= 0;
              imag_value=0;
            end
    12869 : begin
              real_value= 0;
              imag_value=0;
            end
    12870 : begin
              real_value= 0;
              imag_value=0;
            end
    12871 : begin
              real_value= 0;
              imag_value=0;
            end
    12872 : begin
              real_value= 0;
              imag_value=0;
            end
    12873 : begin
              real_value= 0;
              imag_value=0;
            end
    12874 : begin
              real_value= 0;
              imag_value=0;
            end
    12875 : begin
              real_value= 0;
              imag_value=0;
            end
    12876 : begin
              real_value= 0;
              imag_value=0;
            end
    12877 : begin
              real_value= 0;
              imag_value=0;
            end
    12878 : begin
              real_value= 0;
              imag_value=0;
            end
    12879 : begin
              real_value= 0;
              imag_value=0;
            end
    12880 : begin
              real_value= 0;
              imag_value=0;
            end
    12881 : begin
              real_value= 0;
              imag_value=0;
            end
    12882 : begin
              real_value= 0;
              imag_value=0;
            end
    12883 : begin
              real_value= 0;
              imag_value=0;
            end
    12884 : begin
              real_value= 0;
              imag_value=0;
            end
    12885 : begin
              real_value= 0;
              imag_value=0;
            end
    12886 : begin
              real_value= 0;
              imag_value=0;
            end
    12887 : begin
              real_value= 0;
              imag_value=0;
            end
    12888 : begin
              real_value= 0;
              imag_value=0;
            end
    12889 : begin
              real_value= 0;
              imag_value=0;
            end
    12890 : begin
              real_value= 0;
              imag_value=0;
            end
    12891 : begin
              real_value= 0;
              imag_value=0;
            end
    12892 : begin
              real_value= 0;
              imag_value=0;
            end
    12893 : begin
              real_value= 0;
              imag_value=0;
            end
    12894 : begin
              real_value= 0;
              imag_value=0;
            end
    12895 : begin
              real_value= 0;
              imag_value=0;
            end
    12896 : begin
              real_value= 0;
              imag_value=0;
            end
    12897 : begin
              real_value= 0;
              imag_value=0;
            end
    12898 : begin
              real_value= 0;
              imag_value=0;
            end
    12899 : begin
              real_value= 0;
              imag_value=0;
            end
    12900 : begin
              real_value= 0;
              imag_value=0;
            end
    12901 : begin
              real_value= 0;
              imag_value=0;
            end
    12902 : begin
              real_value= 0;
              imag_value=0;
            end
    12903 : begin
              real_value= 0;
              imag_value=0;
            end
    12904 : begin
              real_value= 0;
              imag_value=0;
            end
    12905 : begin
              real_value= 0;
              imag_value=0;
            end
    12906 : begin
              real_value= 0;
              imag_value=0;
            end
    12907 : begin
              real_value= 0;
              imag_value=0;
            end
    12908 : begin
              real_value= 0;
              imag_value=0;
            end
    12909 : begin
              real_value= 0;
              imag_value=0;
            end
    12910 : begin
              real_value= 0;
              imag_value=0;
            end
    12911 : begin
              real_value= 0;
              imag_value=0;
            end
    12912 : begin
              real_value= 0;
              imag_value=0;
            end
    12913 : begin
              real_value= 0;
              imag_value=0;
            end
    12914 : begin
              real_value= 0;
              imag_value=0;
            end
    12915 : begin
              real_value= 0;
              imag_value=0;
            end
    12916 : begin
              real_value= 0;
              imag_value=0;
            end
    12917 : begin
              real_value= 0;
              imag_value=0;
            end
    12918 : begin
              real_value= 0;
              imag_value=0;
            end
    12919 : begin
              real_value= 0;
              imag_value=0;
            end
    12920 : begin
              real_value= 0;
              imag_value=0;
            end
    12921 : begin
              real_value= 0;
              imag_value=0;
            end
    12922 : begin
              real_value= 0;
              imag_value=0;
            end
    12923 : begin
              real_value= 0;
              imag_value=0;
            end
    12924 : begin
              real_value= 0;
              imag_value=0;
            end
    12925 : begin
              real_value= 0;
              imag_value=0;
            end
    12926 : begin
              real_value= 0;
              imag_value=0;
            end
    12927 : begin
              real_value= 0;
              imag_value=0;
            end
    12928 : begin
              real_value= 0;
              imag_value=0;
            end
    12929 : begin
              real_value= 0;
              imag_value=0;
            end
    12930 : begin
              real_value= 0;
              imag_value=0;
            end
    12931 : begin
              real_value= 0;
              imag_value=0;
            end
    12932 : begin
              real_value= 0;
              imag_value=0;
            end
    12933 : begin
              real_value= 0;
              imag_value=0;
            end
    12934 : begin
              real_value= 0;
              imag_value=0;
            end
    12935 : begin
              real_value= 0;
              imag_value=0;
            end
    12936 : begin
              real_value= 0;
              imag_value=0;
            end
    12937 : begin
              real_value= 0;
              imag_value=0;
            end
    12938 : begin
              real_value= 0;
              imag_value=0;
            end
    12939 : begin
              real_value= 0;
              imag_value=0;
            end
    12940 : begin
              real_value= 0;
              imag_value=0;
            end
    12941 : begin
              real_value= 0;
              imag_value=0;
            end
    12942 : begin
              real_value= 0;
              imag_value=0;
            end
    12943 : begin
              real_value= 0;
              imag_value=0;
            end
    12944 : begin
              real_value= 0;
              imag_value=0;
            end
    12945 : begin
              real_value= 0;
              imag_value=0;
            end
    12946 : begin
              real_value= 0;
              imag_value=0;
            end
    12947 : begin
              real_value= 0;
              imag_value=0;
            end
    12948 : begin
              real_value= 0;
              imag_value=0;
            end
    12949 : begin
              real_value= 0;
              imag_value=0;
            end
    12950 : begin
              real_value= 0;
              imag_value=0;
            end
    12951 : begin
              real_value= 0;
              imag_value=0;
            end
    12952 : begin
              real_value= 0;
              imag_value=0;
            end
    12953 : begin
              real_value= 0;
              imag_value=0;
            end
    12954 : begin
              real_value= 0;
              imag_value=0;
            end
    12955 : begin
              real_value= 0;
              imag_value=0;
            end
    12956 : begin
              real_value= 0;
              imag_value=0;
            end
    12957 : begin
              real_value= 0;
              imag_value=0;
            end
    12958 : begin
              real_value= 0;
              imag_value=0;
            end
    12959 : begin
              real_value= 0;
              imag_value=0;
            end
    12960 : begin
              real_value= 0;
              imag_value=0;
            end
    12961 : begin
              real_value= 0;
              imag_value=0;
            end
    12962 : begin
              real_value= 0;
              imag_value=0;
            end
    12963 : begin
              real_value= 0;
              imag_value=0;
            end
    12964 : begin
              real_value= 0;
              imag_value=0;
            end
    12965 : begin
              real_value= 0;
              imag_value=0;
            end
    12966 : begin
              real_value= 0;
              imag_value=0;
            end
    12967 : begin
              real_value= 0;
              imag_value=0;
            end
    12968 : begin
              real_value= 0;
              imag_value=0;
            end
    12969 : begin
              real_value= 0;
              imag_value=0;
            end
    12970 : begin
              real_value= 0;
              imag_value=0;
            end
    12971 : begin
              real_value= 0;
              imag_value=0;
            end
    12972 : begin
              real_value= 0;
              imag_value=0;
            end
    12973 : begin
              real_value= 0;
              imag_value=0;
            end
    12974 : begin
              real_value= 0;
              imag_value=0;
            end
    12975 : begin
              real_value= 0;
              imag_value=0;
            end
    12976 : begin
              real_value= 0;
              imag_value=0;
            end
    12977 : begin
              real_value= 0;
              imag_value=0;
            end
    12978 : begin
              real_value= 0;
              imag_value=0;
            end
    12979 : begin
              real_value= 0;
              imag_value=0;
            end
    12980 : begin
              real_value= 0;
              imag_value=0;
            end
    12981 : begin
              real_value= 0;
              imag_value=0;
            end
    12982 : begin
              real_value= 0;
              imag_value=0;
            end
    12983 : begin
              real_value= 0;
              imag_value=0;
            end
    12984 : begin
              real_value= 0;
              imag_value=0;
            end
    12985 : begin
              real_value= 0;
              imag_value=0;
            end
    12986 : begin
              real_value= 0;
              imag_value=0;
            end
    12987 : begin
              real_value= 0;
              imag_value=0;
            end
    12988 : begin
              real_value= 0;
              imag_value=0;
            end
    12989 : begin
              real_value= 0;
              imag_value=0;
            end
    12990 : begin
              real_value= 0;
              imag_value=0;
            end
    12991 : begin
              real_value= 0;
              imag_value=0;
            end
    12992 : begin
              real_value= 0;
              imag_value=0;
            end
    12993 : begin
              real_value= 0;
              imag_value=0;
            end
    12994 : begin
              real_value= 0;
              imag_value=0;
            end
    12995 : begin
              real_value= 0;
              imag_value=0;
            end
    12996 : begin
              real_value= 0;
              imag_value=0;
            end
    12997 : begin
              real_value= 0;
              imag_value=0;
            end
    12998 : begin
              real_value= 0;
              imag_value=0;
            end
    12999 : begin
              real_value= 0;
              imag_value=0;
            end
    13000 : begin
              real_value= 0;
              imag_value=0;
            end
    13001 : begin
              real_value= 0;
              imag_value=0;
            end
    13002 : begin
              real_value= 0;
              imag_value=0;
            end
    13003 : begin
              real_value= 0;
              imag_value=0;
            end
    13004 : begin
              real_value= 0;
              imag_value=0;
            end
    13005 : begin
              real_value= 0;
              imag_value=0;
            end
    13006 : begin
              real_value= 0;
              imag_value=0;
            end
    13007 : begin
              real_value= 0;
              imag_value=0;
            end
  endcase
end // always @ (*)
   
*/

endmodule   

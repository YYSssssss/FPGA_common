`ifndef _RSP_S1_PREP_DEFINE_SVH_
  `define  _RSP_S1_PREP_DEFINE_SVH_
    `define RSP_S1_PREP_BANK_NUM   14
    `define RSP_S1_PREP_DATA_WIDTH 128
    `define RSP_S1_PREP_ADDR_WIDTH 18
    `define RSP_S1_PREP_STRB_WIDTH 16



`endif

// -------------------------------------------------------------------------- //
// Copyright Jabil Inc.
// -------------------------------------------------------------------------- //
// Name         : Shehanaj Begum                                               //
// Date         : 6/15/20                                                     //
// File         : jb_top_ctrl_test.sv                                                //
// Design       :                                                             //
// Purpose      :                                                             //
// Device       : xczu47dr-fsve1156-2-i-es1                                   //
// -------------------------------------------------------------------------- //

module sensemi_top_ctrl_test #(
    parameter           AXI_ADDR_WIDTH  = 13,
    parameter           AXI_DATA_WIDTH  = 32
)(
    input                       clk,
    input                       srst,
    sensemi_axi4_lite_if.slave       IFP_axi4_lite,
    sensemi_test_ctrl_if.ctrl    IFP_test_ctrl,
    sensemi_test_stat_if.stat    IFP_test_stat 
);

    // ------------------------------------------------------------------ //
    // Register Set: Top Control                                          //
    // ------------------------------------------------------------------ //

    sensemi_axi_regs_if      #(.AXI_ADDR_WIDTH(AXI_ADDR_WIDTH), .AXI_DATA_WIDTH(AXI_DATA_WIDTH)) IFP_axi_rw ();

    sensemi_axi_slave #(
        .AXI_ADDR_WIDTH             (AXI_ADDR_WIDTH),
        .AXI_DATA_WIDTH             (AXI_DATA_WIDTH)
    ) u_axi_slave_top_ctrl (
        .clk                        (clk),                  // i
        .srst                       (srst),                 // i
        .IFP_axi4_lite              (IFP_axi4_lite),     // jb_axi4_lite_if.slave
        .IFP_axi_rw                 (IFP_axi_rw)  // jb_axi_regs_if.master
    );


    sensemi_test_regs u_test_regs (
        .clk                        (clk),                  // i
        .srst                       (srst),                 // i
        .IFP_axi_rw                 (IFP_axi_rw),           // jb_axi_regs_if.slave
        .IFP_test_ctrl              (IFP_test_ctrl),    // mm_regs_top_ctrl_if.ctrl
        .IFP_test_stat              (IFP_test_stat)
    );

    // ------------------------------------------------------------------ //
    // Register Set: ...                                                  //
    // ------------------------------------------------------------------ //

endmodule
 
